*TB DC OTA BUFFERED
.include ../minimal_libs/sky130_libs/sky130_lib.spice
.include ./ota.spice

X1	IN1	IN2	VD	VS	A	OUT ota

CL	OUT	0	4p
*CL	E	0	4p
*CC	D	E	0.88p

Ibias A 0 5.53u

VDD VD 0 1.8
VSS VS 0 -1.8

VIN2 IN2 0 DC 0

*Vin1 com malha aberta
VIN1 IN1 0 DC 1

*Vin1 com malha fechada
*VIN1 R 0 DC 1

*Realimentação
*R1 R IN1 10k
*Rf IN1 E 100k


* cmd 	src	start	stop	step
.dc	VIN1	-1.8	1.8	0.01

.end

.control

run

plot  OUT in1

.endc
