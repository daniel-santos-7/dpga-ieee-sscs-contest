*OTA BUFFERED
.include ../minimal_libs/sky130_libs/sky130_lib.spice

.subckt	ota	in1	in2	vd	vs	ib	out

*label drain   gate    source  bulk   	 model           	length	width   		
XM1      c	in1	b       b	sky130_fd_pr__pfet_01v8  L=1u	W=2.93u
XM2      d	in2	b	b	sky130_fd_pr__pfet_01v8  L=1u	W=2.93u
XM3      c       c	vs	vs	sky130_fd_pr__nfet_01v8  L=1u	W=0.861u
XM4	d	c	vs	vs	sky130_fd_pr__nfet_01v8  L=1u	W=0.861u
XM5	ib	ib	vd	vd	sky130_fd_pr__pfet_01v8  L=1u	W=5.85u
XM6      b	ib	vd	vd	sky130_fd_pr__pfet_01v8  L=1u	W=5.85u
XM7	e	d	vs	vs	sky130_fd_pr__nfet_01v8  L=1u	W=8.61u
XM8	e	ib	vd	vd	sky130_fd_pr__pfet_01v8  L=1u	W=29.3u
XM9	vs	e	out	out	sky130_fd_pr__pfet_01v8  L=1u	W=5.85u
XM10	out	ib	vd	vd	sky130_fd_pr__pfet_01v8  L=1u	W=5.85u

Cc	d	e	0.5p

C0	ib 	b 	2.94fF
C1	ib 	vd 	2.95fF
C2 	d	 b 	430.72fF
C3 	ib 	vs 	3.88fF
C4 	vd 	vs 	2.31fF

.ends
