magic
tech sky130A
magscale 1 2
timestamp 1634766647
<< locali >>
rect 16681 4539 16715 16949
<< viali >>
rect 2421 17221 2455 17255
rect 15485 17221 15519 17255
rect 11713 17153 11747 17187
rect 2605 17017 2639 17051
rect 11529 16949 11563 16983
rect 15761 16949 15795 16983
rect 16681 16949 16715 16983
rect 7757 5185 7791 5219
rect 7849 5185 7883 5219
rect 8125 5185 8159 5219
rect 8769 5185 8803 5219
rect 9597 5185 9631 5219
rect 8033 5049 8067 5083
rect 7573 4981 7607 5015
rect 8585 4981 8619 5015
rect 9689 4981 9723 5015
rect 6929 4641 6963 4675
rect 9045 4641 9079 4675
rect 6653 4573 6687 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 9319 4573 9353 4607
rect 10517 4573 10551 4607
rect 10793 4505 10827 4539
rect 16681 4505 16715 4539
rect 8401 4437 8435 4471
rect 9505 4437 9539 4471
rect 12265 4437 12299 4471
rect 9045 4165 9079 4199
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 12081 4097 12115 4131
rect 12725 4097 12759 4131
rect 12817 4097 12851 4131
rect 13093 4097 13127 4131
rect 6377 4029 6411 4063
rect 6653 4029 6687 4063
rect 11989 4029 12023 4063
rect 8125 3893 8159 3927
rect 10333 3893 10367 3927
rect 11529 3893 11563 3927
rect 12541 3893 12575 3927
rect 13001 3893 13035 3927
rect 8953 3689 8987 3723
rect 5825 3553 5859 3587
rect 10425 3553 10459 3587
rect 10701 3553 10735 3587
rect 11161 3553 11195 3587
rect 11437 3553 11471 3587
rect 5549 3485 5583 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6377 3485 6411 3519
rect 5365 3417 5399 3451
rect 6653 3417 6687 3451
rect 8125 3349 8159 3383
rect 12909 3349 12943 3383
rect 4537 3145 4571 3179
rect 6377 3145 6411 3179
rect 8769 3145 8803 3179
rect 10701 3145 10735 3179
rect 11805 3077 11839 3111
rect 5825 3009 5859 3043
rect 6561 3009 6595 3043
rect 7021 3009 7055 3043
rect 9229 3009 9263 3043
rect 11529 3009 11563 3043
rect 7297 2941 7331 2975
rect 13277 2805 13311 2839
rect 6561 2601 6595 2635
rect 7573 2601 7607 2635
rect 10885 2601 10919 2635
rect 10425 2533 10459 2567
rect 7021 2465 7055 2499
rect 8033 2465 8067 2499
rect 1961 2397 1995 2431
rect 4353 2397 4387 2431
rect 6745 2397 6779 2431
rect 6883 2397 6917 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 9505 2397 9539 2431
rect 10609 2397 10643 2431
rect 10701 2397 10735 2431
rect 10977 2397 11011 2431
rect 11713 2397 11747 2431
rect 12449 2397 12483 2431
rect 14657 2397 14691 2431
rect 15669 2397 15703 2431
rect 1777 2329 1811 2363
rect 4169 2329 4203 2363
rect 5549 2329 5583 2363
rect 5733 2329 5767 2363
rect 11529 2329 11563 2363
rect 12265 2329 12299 2363
rect 14473 2329 14507 2363
rect 15853 2329 15887 2363
rect 9413 2261 9447 2295
<< metal1 >>
rect 1104 17434 16560 17456
rect 1104 17382 6102 17434
rect 6154 17382 6166 17434
rect 6218 17382 6230 17434
rect 6282 17382 6294 17434
rect 6346 17382 6358 17434
rect 6410 17382 11254 17434
rect 11306 17382 11318 17434
rect 11370 17382 11382 17434
rect 11434 17382 11446 17434
rect 11498 17382 11510 17434
rect 11562 17382 16560 17434
rect 1104 17360 16560 17382
rect 2222 17212 2228 17264
rect 2280 17252 2286 17264
rect 2409 17255 2467 17261
rect 2409 17252 2421 17255
rect 2280 17224 2421 17252
rect 2280 17212 2286 17224
rect 2409 17221 2421 17224
rect 2455 17221 2467 17255
rect 15470 17252 15476 17264
rect 15431 17224 15476 17252
rect 2409 17215 2467 17221
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11112 17156 11713 17184
rect 11112 17144 11118 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 2593 17051 2651 17057
rect 2593 17017 2605 17051
rect 2639 17048 2651 17051
rect 7742 17048 7748 17060
rect 2639 17020 7748 17048
rect 2639 17017 2651 17020
rect 2593 17011 2651 17017
rect 7742 17008 7748 17020
rect 7800 17008 7806 17060
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 7892 16952 11529 16980
rect 7892 16940 7898 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 11517 16943 11575 16949
rect 15749 16983 15807 16989
rect 15749 16949 15761 16983
rect 15795 16980 15807 16983
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 15795 16952 16681 16980
rect 15795 16949 15807 16952
rect 15749 16943 15807 16949
rect 16669 16949 16681 16952
rect 16715 16949 16727 16983
rect 16669 16943 16727 16949
rect 1104 16890 16560 16912
rect 1104 16838 3526 16890
rect 3578 16838 3590 16890
rect 3642 16838 3654 16890
rect 3706 16838 3718 16890
rect 3770 16838 3782 16890
rect 3834 16838 8678 16890
rect 8730 16838 8742 16890
rect 8794 16838 8806 16890
rect 8858 16838 8870 16890
rect 8922 16838 8934 16890
rect 8986 16838 13830 16890
rect 13882 16838 13894 16890
rect 13946 16838 13958 16890
rect 14010 16838 14022 16890
rect 14074 16838 14086 16890
rect 14138 16838 16560 16890
rect 1104 16816 16560 16838
rect 1104 16346 16560 16368
rect 1104 16294 6102 16346
rect 6154 16294 6166 16346
rect 6218 16294 6230 16346
rect 6282 16294 6294 16346
rect 6346 16294 6358 16346
rect 6410 16294 11254 16346
rect 11306 16294 11318 16346
rect 11370 16294 11382 16346
rect 11434 16294 11446 16346
rect 11498 16294 11510 16346
rect 11562 16294 16560 16346
rect 1104 16272 16560 16294
rect 1104 15802 16560 15824
rect 1104 15750 3526 15802
rect 3578 15750 3590 15802
rect 3642 15750 3654 15802
rect 3706 15750 3718 15802
rect 3770 15750 3782 15802
rect 3834 15750 8678 15802
rect 8730 15750 8742 15802
rect 8794 15750 8806 15802
rect 8858 15750 8870 15802
rect 8922 15750 8934 15802
rect 8986 15750 13830 15802
rect 13882 15750 13894 15802
rect 13946 15750 13958 15802
rect 14010 15750 14022 15802
rect 14074 15750 14086 15802
rect 14138 15750 16560 15802
rect 1104 15728 16560 15750
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 9030 15348 9036 15360
rect 6696 15320 9036 15348
rect 6696 15308 6702 15320
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 1104 15258 16560 15280
rect 1104 15206 6102 15258
rect 6154 15206 6166 15258
rect 6218 15206 6230 15258
rect 6282 15206 6294 15258
rect 6346 15206 6358 15258
rect 6410 15206 11254 15258
rect 11306 15206 11318 15258
rect 11370 15206 11382 15258
rect 11434 15206 11446 15258
rect 11498 15206 11510 15258
rect 11562 15206 16560 15258
rect 1104 15184 16560 15206
rect 1104 14714 16560 14736
rect 1104 14662 3526 14714
rect 3578 14662 3590 14714
rect 3642 14662 3654 14714
rect 3706 14662 3718 14714
rect 3770 14662 3782 14714
rect 3834 14662 8678 14714
rect 8730 14662 8742 14714
rect 8794 14662 8806 14714
rect 8858 14662 8870 14714
rect 8922 14662 8934 14714
rect 8986 14662 13830 14714
rect 13882 14662 13894 14714
rect 13946 14662 13958 14714
rect 14010 14662 14022 14714
rect 14074 14662 14086 14714
rect 14138 14662 16560 14714
rect 1104 14640 16560 14662
rect 1104 14170 16560 14192
rect 1104 14118 6102 14170
rect 6154 14118 6166 14170
rect 6218 14118 6230 14170
rect 6282 14118 6294 14170
rect 6346 14118 6358 14170
rect 6410 14118 11254 14170
rect 11306 14118 11318 14170
rect 11370 14118 11382 14170
rect 11434 14118 11446 14170
rect 11498 14118 11510 14170
rect 11562 14118 16560 14170
rect 1104 14096 16560 14118
rect 1104 13626 16560 13648
rect 1104 13574 3526 13626
rect 3578 13574 3590 13626
rect 3642 13574 3654 13626
rect 3706 13574 3718 13626
rect 3770 13574 3782 13626
rect 3834 13574 8678 13626
rect 8730 13574 8742 13626
rect 8794 13574 8806 13626
rect 8858 13574 8870 13626
rect 8922 13574 8934 13626
rect 8986 13574 13830 13626
rect 13882 13574 13894 13626
rect 13946 13574 13958 13626
rect 14010 13574 14022 13626
rect 14074 13574 14086 13626
rect 14138 13574 16560 13626
rect 1104 13552 16560 13574
rect 1104 13082 16560 13104
rect 1104 13030 6102 13082
rect 6154 13030 6166 13082
rect 6218 13030 6230 13082
rect 6282 13030 6294 13082
rect 6346 13030 6358 13082
rect 6410 13030 11254 13082
rect 11306 13030 11318 13082
rect 11370 13030 11382 13082
rect 11434 13030 11446 13082
rect 11498 13030 11510 13082
rect 11562 13030 16560 13082
rect 1104 13008 16560 13030
rect 1104 12538 16560 12560
rect 1104 12486 3526 12538
rect 3578 12486 3590 12538
rect 3642 12486 3654 12538
rect 3706 12486 3718 12538
rect 3770 12486 3782 12538
rect 3834 12486 8678 12538
rect 8730 12486 8742 12538
rect 8794 12486 8806 12538
rect 8858 12486 8870 12538
rect 8922 12486 8934 12538
rect 8986 12486 13830 12538
rect 13882 12486 13894 12538
rect 13946 12486 13958 12538
rect 14010 12486 14022 12538
rect 14074 12486 14086 12538
rect 14138 12486 16560 12538
rect 1104 12464 16560 12486
rect 1104 11994 16560 12016
rect 1104 11942 6102 11994
rect 6154 11942 6166 11994
rect 6218 11942 6230 11994
rect 6282 11942 6294 11994
rect 6346 11942 6358 11994
rect 6410 11942 11254 11994
rect 11306 11942 11318 11994
rect 11370 11942 11382 11994
rect 11434 11942 11446 11994
rect 11498 11942 11510 11994
rect 11562 11942 16560 11994
rect 1104 11920 16560 11942
rect 1104 11450 16560 11472
rect 1104 11398 3526 11450
rect 3578 11398 3590 11450
rect 3642 11398 3654 11450
rect 3706 11398 3718 11450
rect 3770 11398 3782 11450
rect 3834 11398 8678 11450
rect 8730 11398 8742 11450
rect 8794 11398 8806 11450
rect 8858 11398 8870 11450
rect 8922 11398 8934 11450
rect 8986 11398 13830 11450
rect 13882 11398 13894 11450
rect 13946 11398 13958 11450
rect 14010 11398 14022 11450
rect 14074 11398 14086 11450
rect 14138 11398 16560 11450
rect 1104 11376 16560 11398
rect 1104 10906 16560 10928
rect 1104 10854 6102 10906
rect 6154 10854 6166 10906
rect 6218 10854 6230 10906
rect 6282 10854 6294 10906
rect 6346 10854 6358 10906
rect 6410 10854 11254 10906
rect 11306 10854 11318 10906
rect 11370 10854 11382 10906
rect 11434 10854 11446 10906
rect 11498 10854 11510 10906
rect 11562 10854 16560 10906
rect 1104 10832 16560 10854
rect 1104 10362 16560 10384
rect 1104 10310 3526 10362
rect 3578 10310 3590 10362
rect 3642 10310 3654 10362
rect 3706 10310 3718 10362
rect 3770 10310 3782 10362
rect 3834 10310 8678 10362
rect 8730 10310 8742 10362
rect 8794 10310 8806 10362
rect 8858 10310 8870 10362
rect 8922 10310 8934 10362
rect 8986 10310 13830 10362
rect 13882 10310 13894 10362
rect 13946 10310 13958 10362
rect 14010 10310 14022 10362
rect 14074 10310 14086 10362
rect 14138 10310 16560 10362
rect 1104 10288 16560 10310
rect 1104 9818 16560 9840
rect 1104 9766 6102 9818
rect 6154 9766 6166 9818
rect 6218 9766 6230 9818
rect 6282 9766 6294 9818
rect 6346 9766 6358 9818
rect 6410 9766 11254 9818
rect 11306 9766 11318 9818
rect 11370 9766 11382 9818
rect 11434 9766 11446 9818
rect 11498 9766 11510 9818
rect 11562 9766 16560 9818
rect 1104 9744 16560 9766
rect 1104 9274 16560 9296
rect 1104 9222 3526 9274
rect 3578 9222 3590 9274
rect 3642 9222 3654 9274
rect 3706 9222 3718 9274
rect 3770 9222 3782 9274
rect 3834 9222 8678 9274
rect 8730 9222 8742 9274
rect 8794 9222 8806 9274
rect 8858 9222 8870 9274
rect 8922 9222 8934 9274
rect 8986 9222 13830 9274
rect 13882 9222 13894 9274
rect 13946 9222 13958 9274
rect 14010 9222 14022 9274
rect 14074 9222 14086 9274
rect 14138 9222 16560 9274
rect 1104 9200 16560 9222
rect 1104 8730 16560 8752
rect 1104 8678 6102 8730
rect 6154 8678 6166 8730
rect 6218 8678 6230 8730
rect 6282 8678 6294 8730
rect 6346 8678 6358 8730
rect 6410 8678 11254 8730
rect 11306 8678 11318 8730
rect 11370 8678 11382 8730
rect 11434 8678 11446 8730
rect 11498 8678 11510 8730
rect 11562 8678 16560 8730
rect 1104 8656 16560 8678
rect 1104 8186 16560 8208
rect 1104 8134 3526 8186
rect 3578 8134 3590 8186
rect 3642 8134 3654 8186
rect 3706 8134 3718 8186
rect 3770 8134 3782 8186
rect 3834 8134 8678 8186
rect 8730 8134 8742 8186
rect 8794 8134 8806 8186
rect 8858 8134 8870 8186
rect 8922 8134 8934 8186
rect 8986 8134 13830 8186
rect 13882 8134 13894 8186
rect 13946 8134 13958 8186
rect 14010 8134 14022 8186
rect 14074 8134 14086 8186
rect 14138 8134 16560 8186
rect 1104 8112 16560 8134
rect 1104 7642 16560 7664
rect 1104 7590 6102 7642
rect 6154 7590 6166 7642
rect 6218 7590 6230 7642
rect 6282 7590 6294 7642
rect 6346 7590 6358 7642
rect 6410 7590 11254 7642
rect 11306 7590 11318 7642
rect 11370 7590 11382 7642
rect 11434 7590 11446 7642
rect 11498 7590 11510 7642
rect 11562 7590 16560 7642
rect 1104 7568 16560 7590
rect 1104 7098 16560 7120
rect 1104 7046 3526 7098
rect 3578 7046 3590 7098
rect 3642 7046 3654 7098
rect 3706 7046 3718 7098
rect 3770 7046 3782 7098
rect 3834 7046 8678 7098
rect 8730 7046 8742 7098
rect 8794 7046 8806 7098
rect 8858 7046 8870 7098
rect 8922 7046 8934 7098
rect 8986 7046 13830 7098
rect 13882 7046 13894 7098
rect 13946 7046 13958 7098
rect 14010 7046 14022 7098
rect 14074 7046 14086 7098
rect 14138 7046 16560 7098
rect 1104 7024 16560 7046
rect 1104 6554 16560 6576
rect 1104 6502 6102 6554
rect 6154 6502 6166 6554
rect 6218 6502 6230 6554
rect 6282 6502 6294 6554
rect 6346 6502 6358 6554
rect 6410 6502 11254 6554
rect 11306 6502 11318 6554
rect 11370 6502 11382 6554
rect 11434 6502 11446 6554
rect 11498 6502 11510 6554
rect 11562 6502 16560 6554
rect 1104 6480 16560 6502
rect 1104 6010 16560 6032
rect 1104 5958 3526 6010
rect 3578 5958 3590 6010
rect 3642 5958 3654 6010
rect 3706 5958 3718 6010
rect 3770 5958 3782 6010
rect 3834 5958 8678 6010
rect 8730 5958 8742 6010
rect 8794 5958 8806 6010
rect 8858 5958 8870 6010
rect 8922 5958 8934 6010
rect 8986 5958 13830 6010
rect 13882 5958 13894 6010
rect 13946 5958 13958 6010
rect 14010 5958 14022 6010
rect 14074 5958 14086 6010
rect 14138 5958 16560 6010
rect 1104 5936 16560 5958
rect 1104 5466 16560 5488
rect 1104 5414 6102 5466
rect 6154 5414 6166 5466
rect 6218 5414 6230 5466
rect 6282 5414 6294 5466
rect 6346 5414 6358 5466
rect 6410 5414 11254 5466
rect 11306 5414 11318 5466
rect 11370 5414 11382 5466
rect 11434 5414 11446 5466
rect 11498 5414 11510 5466
rect 11562 5414 16560 5466
rect 1104 5392 16560 5414
rect 7760 5256 8800 5284
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7760 5225 7788 5256
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7708 5188 7757 5216
rect 7708 5176 7714 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 8113 5219 8171 5225
rect 7892 5188 7937 5216
rect 7892 5176 7898 5188
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8202 5216 8208 5228
rect 8159 5188 8208 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8772 5225 8800 5256
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9585 5219 9643 5225
rect 9585 5216 9597 5219
rect 8803 5188 9597 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9585 5185 9597 5188
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 8021 5083 8079 5089
rect 8021 5080 8033 5083
rect 6880 5052 8033 5080
rect 6880 5040 6886 5052
rect 8021 5049 8033 5052
rect 8067 5049 8079 5083
rect 8021 5043 8079 5049
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 6972 4984 7573 5012
rect 6972 4972 6978 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 8573 5015 8631 5021
rect 8573 4981 8585 5015
rect 8619 5012 8631 5015
rect 9306 5012 9312 5024
rect 8619 4984 9312 5012
rect 8619 4981 8631 4984
rect 8573 4975 8631 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 9674 5012 9680 5024
rect 9635 4984 9680 5012
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 1104 4922 16560 4944
rect 1104 4870 3526 4922
rect 3578 4870 3590 4922
rect 3642 4870 3654 4922
rect 3706 4870 3718 4922
rect 3770 4870 3782 4922
rect 3834 4870 8678 4922
rect 8730 4870 8742 4922
rect 8794 4870 8806 4922
rect 8858 4870 8870 4922
rect 8922 4870 8934 4922
rect 8986 4870 13830 4922
rect 13882 4870 13894 4922
rect 13946 4870 13958 4922
rect 14010 4870 14022 4922
rect 14074 4870 14086 4922
rect 14138 4870 16560 4922
rect 1104 4848 16560 4870
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 9033 4675 9091 4681
rect 6972 4644 7017 4672
rect 6972 4632 6978 4644
rect 9033 4641 9045 4675
rect 9079 4672 9091 4675
rect 9122 4672 9128 4684
rect 9079 4644 9128 4672
rect 9079 4641 9091 4644
rect 9033 4635 9091 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 6454 4564 6460 4616
rect 6512 4604 6518 4616
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 6512 4576 6653 4604
rect 6512 4564 6518 4576
rect 6641 4573 6653 4576
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 8018 4564 8024 4616
rect 8076 4564 8082 4616
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8260 4576 8953 4604
rect 8260 4564 8266 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 8941 4567 8999 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9306 4564 9312 4616
rect 9364 4604 9370 4616
rect 10505 4607 10563 4613
rect 9364 4576 9407 4604
rect 9364 4564 9370 4576
rect 10505 4573 10517 4607
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 6880 4440 8401 4468
rect 6880 4428 6886 4440
rect 8389 4437 8401 4440
rect 8435 4437 8447 4471
rect 8389 4431 8447 4437
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 10410 4468 10416 4480
rect 9539 4440 10416 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10520 4468 10548 4567
rect 10778 4536 10784 4548
rect 10739 4508 10784 4536
rect 10778 4496 10784 4508
rect 10836 4496 10842 4548
rect 12158 4536 12164 4548
rect 12006 4508 12164 4536
rect 12158 4496 12164 4508
rect 12216 4536 12222 4548
rect 16669 4539 16727 4545
rect 16669 4536 16681 4539
rect 12216 4508 16681 4536
rect 12216 4496 12222 4508
rect 16669 4505 16681 4508
rect 16715 4505 16727 4539
rect 16669 4499 16727 4505
rect 10686 4468 10692 4480
rect 10520 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 12253 4471 12311 4477
rect 12253 4437 12265 4471
rect 12299 4468 12311 4471
rect 12342 4468 12348 4480
rect 12299 4440 12348 4468
rect 12299 4437 12311 4440
rect 12253 4431 12311 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 1104 4378 16560 4400
rect 1104 4326 6102 4378
rect 6154 4326 6166 4378
rect 6218 4326 6230 4378
rect 6282 4326 6294 4378
rect 6346 4326 6358 4378
rect 6410 4326 11254 4378
rect 11306 4326 11318 4378
rect 11370 4326 11382 4378
rect 11434 4326 11446 4378
rect 11498 4326 11510 4378
rect 11562 4326 16560 4378
rect 1104 4304 16560 4326
rect 8018 4196 8024 4208
rect 7866 4168 8024 4196
rect 8018 4156 8024 4168
rect 8076 4156 8082 4208
rect 9030 4196 9036 4208
rect 8991 4168 9036 4196
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 9364 4168 12848 4196
rect 9364 4156 9370 4168
rect 11716 4137 11744 4168
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12069 4131 12127 4137
rect 11848 4100 11893 4128
rect 11848 4088 11854 4100
rect 12069 4097 12081 4131
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 6362 4060 6368 4072
rect 6323 4032 6368 4060
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 6638 4060 6644 4072
rect 6599 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 9674 4060 9680 4072
rect 6788 4032 9680 4060
rect 6788 4020 6794 4032
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 10870 4060 10876 4072
rect 9732 4032 10876 4060
rect 9732 4020 9738 4032
rect 10870 4020 10876 4032
rect 10928 4060 10934 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 10928 4032 11989 4060
rect 10928 4020 10934 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 12084 4060 12112 4091
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12820 4137 12848 4168
rect 12713 4131 12771 4137
rect 12713 4128 12725 4131
rect 12400 4100 12725 4128
rect 12400 4088 12406 4100
rect 12713 4097 12725 4100
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4097 12863 4131
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12805 4091 12863 4097
rect 13004 4100 13093 4128
rect 12434 4060 12440 4072
rect 12084 4032 12440 4060
rect 11977 4023 12035 4029
rect 11992 3992 12020 4023
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 13004 3992 13032 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 11992 3964 13032 3992
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11480 3896 11529 3924
rect 11480 3884 11486 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12124 3896 12541 3924
rect 12124 3884 12130 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12529 3887 12587 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 1104 3834 16560 3856
rect 1104 3782 3526 3834
rect 3578 3782 3590 3834
rect 3642 3782 3654 3834
rect 3706 3782 3718 3834
rect 3770 3782 3782 3834
rect 3834 3782 8678 3834
rect 8730 3782 8742 3834
rect 8794 3782 8806 3834
rect 8858 3782 8870 3834
rect 8922 3782 8934 3834
rect 8986 3782 13830 3834
rect 13882 3782 13894 3834
rect 13946 3782 13958 3834
rect 14010 3782 14022 3834
rect 14074 3782 14086 3834
rect 14138 3782 16560 3834
rect 1104 3760 16560 3782
rect 7006 3720 7012 3732
rect 5644 3692 7012 3720
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 5644 3525 5672 3692
rect 7006 3680 7012 3692
rect 7064 3720 7070 3732
rect 8110 3720 8116 3732
rect 7064 3692 8116 3720
rect 7064 3680 7070 3692
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9122 3720 9128 3732
rect 8987 3692 9128 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9122 3680 9128 3692
rect 9180 3720 9186 3732
rect 11790 3720 11796 3732
rect 9180 3692 11796 3720
rect 9180 3680 9186 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 7926 3584 7932 3596
rect 5859 3556 7932 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 10410 3584 10416 3596
rect 10371 3556 10416 3584
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3584 10750 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10744 3556 11161 3584
rect 10744 3544 10750 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11422 3584 11428 3596
rect 11383 3556 11428 3584
rect 11149 3547 11207 3553
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 5629 3479 5687 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6362 3516 6368 3528
rect 6052 3488 6368 3516
rect 6052 3476 6058 3488
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 6641 3451 6699 3457
rect 6641 3448 6653 3451
rect 5399 3420 6653 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6641 3417 6653 3420
rect 6687 3417 6699 3451
rect 8018 3448 8024 3460
rect 7866 3420 8024 3448
rect 6641 3411 6699 3417
rect 8018 3408 8024 3420
rect 8076 3448 8082 3460
rect 8076 3420 8248 3448
rect 8076 3408 8082 3420
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 6546 3380 6552 3392
rect 5592 3352 6552 3380
rect 5592 3340 5598 3352
rect 6546 3340 6552 3352
rect 6604 3380 6610 3392
rect 7650 3380 7656 3392
rect 6604 3352 7656 3380
rect 6604 3340 6610 3352
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 7984 3352 8125 3380
rect 7984 3340 7990 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8220 3380 8248 3420
rect 9968 3380 9996 3434
rect 12158 3408 12164 3460
rect 12216 3408 12222 3460
rect 12176 3380 12204 3408
rect 8220 3352 12204 3380
rect 8113 3343 8171 3349
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12897 3383 12955 3389
rect 12897 3380 12909 3383
rect 12492 3352 12909 3380
rect 12492 3340 12498 3352
rect 12897 3349 12909 3352
rect 12943 3349 12955 3383
rect 12897 3343 12955 3349
rect 1104 3290 16560 3312
rect 1104 3238 6102 3290
rect 6154 3238 6166 3290
rect 6218 3238 6230 3290
rect 6282 3238 6294 3290
rect 6346 3238 6358 3290
rect 6410 3238 11254 3290
rect 11306 3238 11318 3290
rect 11370 3238 11382 3290
rect 11434 3238 11446 3290
rect 11498 3238 11510 3290
rect 11562 3238 16560 3290
rect 1104 3216 16560 3238
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 4540 3108 4568 3139
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5960 3148 6377 3176
rect 5960 3136 5966 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9214 3176 9220 3188
rect 8803 3148 9220 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 10686 3176 10692 3188
rect 10647 3148 10692 3176
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 12158 3136 12164 3188
rect 12216 3136 12222 3188
rect 5994 3108 6000 3120
rect 4540 3080 6000 3108
rect 5994 3068 6000 3080
rect 6052 3108 6058 3120
rect 6052 3080 6914 3108
rect 6052 3068 6058 3080
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 6730 3040 6736 3052
rect 6595 3012 6736 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 5828 2904 5856 3003
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 6886 3040 6914 3080
rect 8018 3068 8024 3120
rect 8076 3068 8082 3120
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6886 3012 7021 3040
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3040 9275 3043
rect 10318 3040 10324 3052
rect 9263 3012 10324 3040
rect 9263 3009 9275 3012
rect 9217 3003 9275 3009
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 5828 2876 7144 2904
rect 5902 2796 5908 2848
rect 5960 2836 5966 2848
rect 6914 2836 6920 2848
rect 5960 2808 6920 2836
rect 5960 2796 5966 2808
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7116 2836 7144 2876
rect 9232 2836 9260 3003
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10704 3040 10732 3136
rect 11793 3111 11851 3117
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 12066 3108 12072 3120
rect 11839 3080 12072 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 12176 3108 12204 3136
rect 12176 3080 12282 3108
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 10704 3012 11529 3040
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 7116 2808 9260 2836
rect 12986 2796 12992 2848
rect 13044 2836 13050 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 13044 2808 13277 2836
rect 13044 2796 13050 2808
rect 13265 2805 13277 2808
rect 13311 2836 13323 2839
rect 15654 2836 15660 2848
rect 13311 2808 15660 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 1104 2746 16560 2768
rect 1104 2694 3526 2746
rect 3578 2694 3590 2746
rect 3642 2694 3654 2746
rect 3706 2694 3718 2746
rect 3770 2694 3782 2746
rect 3834 2694 8678 2746
rect 8730 2694 8742 2746
rect 8794 2694 8806 2746
rect 8858 2694 8870 2746
rect 8922 2694 8934 2746
rect 8986 2694 13830 2746
rect 13882 2694 13894 2746
rect 13946 2694 13958 2746
rect 14010 2694 14022 2746
rect 14074 2694 14086 2746
rect 14138 2694 16560 2746
rect 1104 2672 16560 2694
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6638 2632 6644 2644
rect 6595 2604 6644 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7340 2604 7573 2632
rect 7340 2592 7346 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 10870 2632 10876 2644
rect 10831 2604 10876 2632
rect 7561 2595 7619 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 6822 2564 6828 2576
rect 1964 2536 6828 2564
rect 1964 2437 1992 2536
rect 6822 2524 6828 2536
rect 6880 2564 6886 2576
rect 9306 2564 9312 2576
rect 6880 2524 6914 2564
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4387 2400 6500 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 1118 2320 1124 2372
rect 1176 2360 1182 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1176 2332 1777 2360
rect 1176 2320 1182 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 3326 2320 3332 2372
rect 3384 2360 3390 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3384 2332 4169 2360
rect 3384 2320 3390 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 5534 2360 5540 2372
rect 5495 2332 5540 2360
rect 4157 2323 4215 2329
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 5721 2363 5779 2369
rect 5721 2329 5733 2363
rect 5767 2329 5779 2363
rect 6472 2360 6500 2400
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 6886 2437 6914 2524
rect 7760 2536 9312 2564
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7064 2468 7157 2496
rect 7064 2456 7070 2468
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6604 2400 6745 2428
rect 6604 2388 6610 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6871 2431 6929 2437
rect 6871 2397 6883 2431
rect 6917 2397 6929 2431
rect 6871 2391 6929 2397
rect 7024 2360 7052 2456
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7760 2437 7788 2536
rect 9306 2524 9312 2536
rect 9364 2564 9370 2576
rect 10413 2567 10471 2573
rect 9364 2536 10364 2564
rect 9364 2524 9370 2536
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 9214 2496 9220 2508
rect 8067 2468 9220 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 9214 2456 9220 2468
rect 9272 2496 9278 2508
rect 10336 2496 10364 2536
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 10778 2564 10784 2576
rect 10459 2536 10784 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 12342 2564 12348 2576
rect 10980 2536 12348 2564
rect 9272 2468 9536 2496
rect 10336 2468 10732 2496
rect 9272 2456 9278 2468
rect 7745 2431 7803 2437
rect 7156 2400 7201 2428
rect 7156 2388 7162 2400
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8113 2431 8171 2437
rect 7892 2400 7937 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 8202 2428 8208 2440
rect 8159 2400 8208 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 6472 2332 7052 2360
rect 7116 2360 7144 2388
rect 8128 2360 8156 2391
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 9508 2437 9536 2468
rect 10704 2437 10732 2468
rect 10980 2437 11008 2536
rect 12342 2524 12348 2536
rect 12400 2564 12406 2576
rect 12400 2536 14688 2564
rect 12400 2524 12406 2536
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 11790 2428 11796 2440
rect 11747 2400 11796 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 7116 2332 8156 2360
rect 5721 2323 5779 2329
rect 5736 2292 5764 2323
rect 7650 2292 7656 2304
rect 5736 2264 7656 2292
rect 7650 2252 7656 2264
rect 7708 2252 7714 2304
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 7800 2264 9413 2292
rect 7800 2252 7806 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 10612 2292 10640 2391
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12434 2388 12440 2440
rect 12492 2428 12498 2440
rect 14660 2437 14688 2536
rect 14645 2431 14703 2437
rect 12492 2400 12537 2428
rect 12492 2388 12498 2400
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 15654 2428 15660 2440
rect 15615 2400 15660 2428
rect 14645 2391 14703 2397
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 10778 2320 10784 2372
rect 10836 2360 10842 2372
rect 11517 2363 11575 2369
rect 11517 2360 11529 2363
rect 10836 2332 11529 2360
rect 10836 2320 10842 2332
rect 11517 2329 11529 2332
rect 11563 2329 11575 2363
rect 11517 2323 11575 2329
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 12253 2363 12311 2369
rect 12253 2360 12265 2363
rect 12216 2332 12265 2360
rect 12216 2320 12222 2332
rect 12253 2329 12265 2332
rect 12299 2329 12311 2363
rect 12253 2323 12311 2329
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 14424 2332 14473 2360
rect 14424 2320 14430 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 15841 2363 15899 2369
rect 15841 2329 15853 2363
rect 15887 2360 15899 2363
rect 16574 2360 16580 2372
rect 15887 2332 16580 2360
rect 15887 2329 15899 2332
rect 15841 2323 15899 2329
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 12434 2292 12440 2304
rect 10612 2264 12440 2292
rect 9401 2255 9459 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 1104 2202 16560 2224
rect 1104 2150 6102 2202
rect 6154 2150 6166 2202
rect 6218 2150 6230 2202
rect 6282 2150 6294 2202
rect 6346 2150 6358 2202
rect 6410 2150 11254 2202
rect 11306 2150 11318 2202
rect 11370 2150 11382 2202
rect 11434 2150 11446 2202
rect 11498 2150 11510 2202
rect 11562 2150 16560 2202
rect 1104 2128 16560 2150
<< via1 >>
rect 6102 17382 6154 17434
rect 6166 17382 6218 17434
rect 6230 17382 6282 17434
rect 6294 17382 6346 17434
rect 6358 17382 6410 17434
rect 11254 17382 11306 17434
rect 11318 17382 11370 17434
rect 11382 17382 11434 17434
rect 11446 17382 11498 17434
rect 11510 17382 11562 17434
rect 2228 17212 2280 17264
rect 15476 17255 15528 17264
rect 15476 17221 15485 17255
rect 15485 17221 15519 17255
rect 15519 17221 15528 17255
rect 15476 17212 15528 17221
rect 11060 17144 11112 17196
rect 7748 17008 7800 17060
rect 7840 16940 7892 16992
rect 3526 16838 3578 16890
rect 3590 16838 3642 16890
rect 3654 16838 3706 16890
rect 3718 16838 3770 16890
rect 3782 16838 3834 16890
rect 8678 16838 8730 16890
rect 8742 16838 8794 16890
rect 8806 16838 8858 16890
rect 8870 16838 8922 16890
rect 8934 16838 8986 16890
rect 13830 16838 13882 16890
rect 13894 16838 13946 16890
rect 13958 16838 14010 16890
rect 14022 16838 14074 16890
rect 14086 16838 14138 16890
rect 6102 16294 6154 16346
rect 6166 16294 6218 16346
rect 6230 16294 6282 16346
rect 6294 16294 6346 16346
rect 6358 16294 6410 16346
rect 11254 16294 11306 16346
rect 11318 16294 11370 16346
rect 11382 16294 11434 16346
rect 11446 16294 11498 16346
rect 11510 16294 11562 16346
rect 3526 15750 3578 15802
rect 3590 15750 3642 15802
rect 3654 15750 3706 15802
rect 3718 15750 3770 15802
rect 3782 15750 3834 15802
rect 8678 15750 8730 15802
rect 8742 15750 8794 15802
rect 8806 15750 8858 15802
rect 8870 15750 8922 15802
rect 8934 15750 8986 15802
rect 13830 15750 13882 15802
rect 13894 15750 13946 15802
rect 13958 15750 14010 15802
rect 14022 15750 14074 15802
rect 14086 15750 14138 15802
rect 6644 15308 6696 15360
rect 9036 15308 9088 15360
rect 6102 15206 6154 15258
rect 6166 15206 6218 15258
rect 6230 15206 6282 15258
rect 6294 15206 6346 15258
rect 6358 15206 6410 15258
rect 11254 15206 11306 15258
rect 11318 15206 11370 15258
rect 11382 15206 11434 15258
rect 11446 15206 11498 15258
rect 11510 15206 11562 15258
rect 3526 14662 3578 14714
rect 3590 14662 3642 14714
rect 3654 14662 3706 14714
rect 3718 14662 3770 14714
rect 3782 14662 3834 14714
rect 8678 14662 8730 14714
rect 8742 14662 8794 14714
rect 8806 14662 8858 14714
rect 8870 14662 8922 14714
rect 8934 14662 8986 14714
rect 13830 14662 13882 14714
rect 13894 14662 13946 14714
rect 13958 14662 14010 14714
rect 14022 14662 14074 14714
rect 14086 14662 14138 14714
rect 6102 14118 6154 14170
rect 6166 14118 6218 14170
rect 6230 14118 6282 14170
rect 6294 14118 6346 14170
rect 6358 14118 6410 14170
rect 11254 14118 11306 14170
rect 11318 14118 11370 14170
rect 11382 14118 11434 14170
rect 11446 14118 11498 14170
rect 11510 14118 11562 14170
rect 3526 13574 3578 13626
rect 3590 13574 3642 13626
rect 3654 13574 3706 13626
rect 3718 13574 3770 13626
rect 3782 13574 3834 13626
rect 8678 13574 8730 13626
rect 8742 13574 8794 13626
rect 8806 13574 8858 13626
rect 8870 13574 8922 13626
rect 8934 13574 8986 13626
rect 13830 13574 13882 13626
rect 13894 13574 13946 13626
rect 13958 13574 14010 13626
rect 14022 13574 14074 13626
rect 14086 13574 14138 13626
rect 6102 13030 6154 13082
rect 6166 13030 6218 13082
rect 6230 13030 6282 13082
rect 6294 13030 6346 13082
rect 6358 13030 6410 13082
rect 11254 13030 11306 13082
rect 11318 13030 11370 13082
rect 11382 13030 11434 13082
rect 11446 13030 11498 13082
rect 11510 13030 11562 13082
rect 3526 12486 3578 12538
rect 3590 12486 3642 12538
rect 3654 12486 3706 12538
rect 3718 12486 3770 12538
rect 3782 12486 3834 12538
rect 8678 12486 8730 12538
rect 8742 12486 8794 12538
rect 8806 12486 8858 12538
rect 8870 12486 8922 12538
rect 8934 12486 8986 12538
rect 13830 12486 13882 12538
rect 13894 12486 13946 12538
rect 13958 12486 14010 12538
rect 14022 12486 14074 12538
rect 14086 12486 14138 12538
rect 6102 11942 6154 11994
rect 6166 11942 6218 11994
rect 6230 11942 6282 11994
rect 6294 11942 6346 11994
rect 6358 11942 6410 11994
rect 11254 11942 11306 11994
rect 11318 11942 11370 11994
rect 11382 11942 11434 11994
rect 11446 11942 11498 11994
rect 11510 11942 11562 11994
rect 3526 11398 3578 11450
rect 3590 11398 3642 11450
rect 3654 11398 3706 11450
rect 3718 11398 3770 11450
rect 3782 11398 3834 11450
rect 8678 11398 8730 11450
rect 8742 11398 8794 11450
rect 8806 11398 8858 11450
rect 8870 11398 8922 11450
rect 8934 11398 8986 11450
rect 13830 11398 13882 11450
rect 13894 11398 13946 11450
rect 13958 11398 14010 11450
rect 14022 11398 14074 11450
rect 14086 11398 14138 11450
rect 6102 10854 6154 10906
rect 6166 10854 6218 10906
rect 6230 10854 6282 10906
rect 6294 10854 6346 10906
rect 6358 10854 6410 10906
rect 11254 10854 11306 10906
rect 11318 10854 11370 10906
rect 11382 10854 11434 10906
rect 11446 10854 11498 10906
rect 11510 10854 11562 10906
rect 3526 10310 3578 10362
rect 3590 10310 3642 10362
rect 3654 10310 3706 10362
rect 3718 10310 3770 10362
rect 3782 10310 3834 10362
rect 8678 10310 8730 10362
rect 8742 10310 8794 10362
rect 8806 10310 8858 10362
rect 8870 10310 8922 10362
rect 8934 10310 8986 10362
rect 13830 10310 13882 10362
rect 13894 10310 13946 10362
rect 13958 10310 14010 10362
rect 14022 10310 14074 10362
rect 14086 10310 14138 10362
rect 6102 9766 6154 9818
rect 6166 9766 6218 9818
rect 6230 9766 6282 9818
rect 6294 9766 6346 9818
rect 6358 9766 6410 9818
rect 11254 9766 11306 9818
rect 11318 9766 11370 9818
rect 11382 9766 11434 9818
rect 11446 9766 11498 9818
rect 11510 9766 11562 9818
rect 3526 9222 3578 9274
rect 3590 9222 3642 9274
rect 3654 9222 3706 9274
rect 3718 9222 3770 9274
rect 3782 9222 3834 9274
rect 8678 9222 8730 9274
rect 8742 9222 8794 9274
rect 8806 9222 8858 9274
rect 8870 9222 8922 9274
rect 8934 9222 8986 9274
rect 13830 9222 13882 9274
rect 13894 9222 13946 9274
rect 13958 9222 14010 9274
rect 14022 9222 14074 9274
rect 14086 9222 14138 9274
rect 6102 8678 6154 8730
rect 6166 8678 6218 8730
rect 6230 8678 6282 8730
rect 6294 8678 6346 8730
rect 6358 8678 6410 8730
rect 11254 8678 11306 8730
rect 11318 8678 11370 8730
rect 11382 8678 11434 8730
rect 11446 8678 11498 8730
rect 11510 8678 11562 8730
rect 3526 8134 3578 8186
rect 3590 8134 3642 8186
rect 3654 8134 3706 8186
rect 3718 8134 3770 8186
rect 3782 8134 3834 8186
rect 8678 8134 8730 8186
rect 8742 8134 8794 8186
rect 8806 8134 8858 8186
rect 8870 8134 8922 8186
rect 8934 8134 8986 8186
rect 13830 8134 13882 8186
rect 13894 8134 13946 8186
rect 13958 8134 14010 8186
rect 14022 8134 14074 8186
rect 14086 8134 14138 8186
rect 6102 7590 6154 7642
rect 6166 7590 6218 7642
rect 6230 7590 6282 7642
rect 6294 7590 6346 7642
rect 6358 7590 6410 7642
rect 11254 7590 11306 7642
rect 11318 7590 11370 7642
rect 11382 7590 11434 7642
rect 11446 7590 11498 7642
rect 11510 7590 11562 7642
rect 3526 7046 3578 7098
rect 3590 7046 3642 7098
rect 3654 7046 3706 7098
rect 3718 7046 3770 7098
rect 3782 7046 3834 7098
rect 8678 7046 8730 7098
rect 8742 7046 8794 7098
rect 8806 7046 8858 7098
rect 8870 7046 8922 7098
rect 8934 7046 8986 7098
rect 13830 7046 13882 7098
rect 13894 7046 13946 7098
rect 13958 7046 14010 7098
rect 14022 7046 14074 7098
rect 14086 7046 14138 7098
rect 6102 6502 6154 6554
rect 6166 6502 6218 6554
rect 6230 6502 6282 6554
rect 6294 6502 6346 6554
rect 6358 6502 6410 6554
rect 11254 6502 11306 6554
rect 11318 6502 11370 6554
rect 11382 6502 11434 6554
rect 11446 6502 11498 6554
rect 11510 6502 11562 6554
rect 3526 5958 3578 6010
rect 3590 5958 3642 6010
rect 3654 5958 3706 6010
rect 3718 5958 3770 6010
rect 3782 5958 3834 6010
rect 8678 5958 8730 6010
rect 8742 5958 8794 6010
rect 8806 5958 8858 6010
rect 8870 5958 8922 6010
rect 8934 5958 8986 6010
rect 13830 5958 13882 6010
rect 13894 5958 13946 6010
rect 13958 5958 14010 6010
rect 14022 5958 14074 6010
rect 14086 5958 14138 6010
rect 6102 5414 6154 5466
rect 6166 5414 6218 5466
rect 6230 5414 6282 5466
rect 6294 5414 6346 5466
rect 6358 5414 6410 5466
rect 11254 5414 11306 5466
rect 11318 5414 11370 5466
rect 11382 5414 11434 5466
rect 11446 5414 11498 5466
rect 11510 5414 11562 5466
rect 7656 5176 7708 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8208 5176 8260 5228
rect 6828 5040 6880 5092
rect 6920 4972 6972 5024
rect 9312 4972 9364 5024
rect 9680 5015 9732 5024
rect 9680 4981 9689 5015
rect 9689 4981 9723 5015
rect 9723 4981 9732 5015
rect 9680 4972 9732 4981
rect 3526 4870 3578 4922
rect 3590 4870 3642 4922
rect 3654 4870 3706 4922
rect 3718 4870 3770 4922
rect 3782 4870 3834 4922
rect 8678 4870 8730 4922
rect 8742 4870 8794 4922
rect 8806 4870 8858 4922
rect 8870 4870 8922 4922
rect 8934 4870 8986 4922
rect 13830 4870 13882 4922
rect 13894 4870 13946 4922
rect 13958 4870 14010 4922
rect 14022 4870 14074 4922
rect 14086 4870 14138 4922
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 9128 4632 9180 4684
rect 6460 4564 6512 4616
rect 8024 4564 8076 4616
rect 8208 4564 8260 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9312 4607 9364 4616
rect 9312 4573 9319 4607
rect 9319 4573 9353 4607
rect 9353 4573 9364 4607
rect 9312 4564 9364 4573
rect 6828 4428 6880 4480
rect 10416 4428 10468 4480
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 12164 4496 12216 4548
rect 10692 4428 10744 4480
rect 12348 4428 12400 4480
rect 6102 4326 6154 4378
rect 6166 4326 6218 4378
rect 6230 4326 6282 4378
rect 6294 4326 6346 4378
rect 6358 4326 6410 4378
rect 11254 4326 11306 4378
rect 11318 4326 11370 4378
rect 11382 4326 11434 4378
rect 11446 4326 11498 4378
rect 11510 4326 11562 4378
rect 8024 4156 8076 4208
rect 9036 4199 9088 4208
rect 9036 4165 9045 4199
rect 9045 4165 9079 4199
rect 9079 4165 9088 4199
rect 9036 4156 9088 4165
rect 9312 4156 9364 4208
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 6368 4063 6420 4072
rect 6368 4029 6377 4063
rect 6377 4029 6411 4063
rect 6411 4029 6420 4063
rect 6368 4020 6420 4029
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 6736 4020 6788 4072
rect 9680 4020 9732 4072
rect 10876 4020 10928 4072
rect 12348 4088 12400 4140
rect 12440 4020 12492 4072
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11428 3884 11480 3936
rect 12072 3884 12124 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 3526 3782 3578 3834
rect 3590 3782 3642 3834
rect 3654 3782 3706 3834
rect 3718 3782 3770 3834
rect 3782 3782 3834 3834
rect 8678 3782 8730 3834
rect 8742 3782 8794 3834
rect 8806 3782 8858 3834
rect 8870 3782 8922 3834
rect 8934 3782 8986 3834
rect 13830 3782 13882 3834
rect 13894 3782 13946 3834
rect 13958 3782 14010 3834
rect 14022 3782 14074 3834
rect 14086 3782 14138 3834
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7012 3680 7064 3732
rect 8116 3680 8168 3732
rect 9128 3680 9180 3732
rect 11796 3680 11848 3732
rect 7932 3544 7984 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 11428 3587 11480 3596
rect 11428 3553 11437 3587
rect 11437 3553 11471 3587
rect 11471 3553 11480 3587
rect 11428 3544 11480 3553
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6000 3476 6052 3528
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 8024 3408 8076 3460
rect 5540 3340 5592 3392
rect 6552 3340 6604 3392
rect 7656 3340 7708 3392
rect 7932 3340 7984 3392
rect 12164 3408 12216 3460
rect 12440 3340 12492 3392
rect 6102 3238 6154 3290
rect 6166 3238 6218 3290
rect 6230 3238 6282 3290
rect 6294 3238 6346 3290
rect 6358 3238 6410 3290
rect 11254 3238 11306 3290
rect 11318 3238 11370 3290
rect 11382 3238 11434 3290
rect 11446 3238 11498 3290
rect 11510 3238 11562 3290
rect 5908 3136 5960 3188
rect 9220 3136 9272 3188
rect 10692 3179 10744 3188
rect 10692 3145 10701 3179
rect 10701 3145 10735 3179
rect 10735 3145 10744 3179
rect 10692 3136 10744 3145
rect 12164 3136 12216 3188
rect 6000 3068 6052 3120
rect 6736 3000 6788 3052
rect 8024 3068 8076 3120
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 5908 2796 5960 2848
rect 6920 2796 6972 2848
rect 10324 3000 10376 3052
rect 12072 3068 12124 3120
rect 12992 2796 13044 2848
rect 15660 2796 15712 2848
rect 3526 2694 3578 2746
rect 3590 2694 3642 2746
rect 3654 2694 3706 2746
rect 3718 2694 3770 2746
rect 3782 2694 3834 2746
rect 8678 2694 8730 2746
rect 8742 2694 8794 2746
rect 8806 2694 8858 2746
rect 8870 2694 8922 2746
rect 8934 2694 8986 2746
rect 13830 2694 13882 2746
rect 13894 2694 13946 2746
rect 13958 2694 14010 2746
rect 14022 2694 14074 2746
rect 14086 2694 14138 2746
rect 6644 2592 6696 2644
rect 7288 2592 7340 2644
rect 10876 2635 10928 2644
rect 10876 2601 10885 2635
rect 10885 2601 10919 2635
rect 10919 2601 10928 2635
rect 10876 2592 10928 2601
rect 6828 2524 6880 2576
rect 1124 2320 1176 2372
rect 3332 2320 3384 2372
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 6552 2388 6604 2440
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 9312 2524 9364 2576
rect 9220 2456 9272 2508
rect 10784 2524 10836 2576
rect 7104 2388 7156 2397
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8208 2388 8260 2440
rect 12348 2524 12400 2576
rect 7656 2252 7708 2304
rect 7748 2252 7800 2304
rect 11796 2388 11848 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 10784 2320 10836 2372
rect 12164 2320 12216 2372
rect 14372 2320 14424 2372
rect 16580 2320 16632 2372
rect 12440 2252 12492 2304
rect 6102 2150 6154 2202
rect 6166 2150 6218 2202
rect 6230 2150 6282 2202
rect 6294 2150 6346 2202
rect 6358 2150 6410 2202
rect 11254 2150 11306 2202
rect 11318 2150 11370 2202
rect 11382 2150 11434 2202
rect 11446 2150 11498 2202
rect 11510 2150 11562 2202
<< metal2 >>
rect 2226 19084 2282 19884
rect 6642 19084 6698 19884
rect 11058 19084 11114 19884
rect 15474 19084 15530 19884
rect 2240 17270 2268 19084
rect 6102 17436 6410 17456
rect 6102 17434 6108 17436
rect 6164 17434 6188 17436
rect 6244 17434 6268 17436
rect 6324 17434 6348 17436
rect 6404 17434 6410 17436
rect 6164 17382 6166 17434
rect 6346 17382 6348 17434
rect 6102 17380 6108 17382
rect 6164 17380 6188 17382
rect 6244 17380 6268 17382
rect 6324 17380 6348 17382
rect 6404 17380 6410 17382
rect 6102 17360 6410 17380
rect 2228 17264 2280 17270
rect 2228 17206 2280 17212
rect 3526 16892 3834 16912
rect 3526 16890 3532 16892
rect 3588 16890 3612 16892
rect 3668 16890 3692 16892
rect 3748 16890 3772 16892
rect 3828 16890 3834 16892
rect 3588 16838 3590 16890
rect 3770 16838 3772 16890
rect 3526 16836 3532 16838
rect 3588 16836 3612 16838
rect 3668 16836 3692 16838
rect 3748 16836 3772 16838
rect 3828 16836 3834 16838
rect 3526 16816 3834 16836
rect 6102 16348 6410 16368
rect 6102 16346 6108 16348
rect 6164 16346 6188 16348
rect 6244 16346 6268 16348
rect 6324 16346 6348 16348
rect 6404 16346 6410 16348
rect 6164 16294 6166 16346
rect 6346 16294 6348 16346
rect 6102 16292 6108 16294
rect 6164 16292 6188 16294
rect 6244 16292 6268 16294
rect 6324 16292 6348 16294
rect 6404 16292 6410 16294
rect 6102 16272 6410 16292
rect 3526 15804 3834 15824
rect 3526 15802 3532 15804
rect 3588 15802 3612 15804
rect 3668 15802 3692 15804
rect 3748 15802 3772 15804
rect 3828 15802 3834 15804
rect 3588 15750 3590 15802
rect 3770 15750 3772 15802
rect 3526 15748 3532 15750
rect 3588 15748 3612 15750
rect 3668 15748 3692 15750
rect 3748 15748 3772 15750
rect 3828 15748 3834 15750
rect 3526 15728 3834 15748
rect 6656 15366 6684 19084
rect 11072 17202 11100 19084
rect 11254 17436 11562 17456
rect 11254 17434 11260 17436
rect 11316 17434 11340 17436
rect 11396 17434 11420 17436
rect 11476 17434 11500 17436
rect 11556 17434 11562 17436
rect 11316 17382 11318 17434
rect 11498 17382 11500 17434
rect 11254 17380 11260 17382
rect 11316 17380 11340 17382
rect 11396 17380 11420 17382
rect 11476 17380 11500 17382
rect 11556 17380 11562 17382
rect 11254 17360 11562 17380
rect 15488 17270 15516 19084
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6102 15260 6410 15280
rect 6102 15258 6108 15260
rect 6164 15258 6188 15260
rect 6244 15258 6268 15260
rect 6324 15258 6348 15260
rect 6404 15258 6410 15260
rect 6164 15206 6166 15258
rect 6346 15206 6348 15258
rect 6102 15204 6108 15206
rect 6164 15204 6188 15206
rect 6244 15204 6268 15206
rect 6324 15204 6348 15206
rect 6404 15204 6410 15206
rect 6102 15184 6410 15204
rect 3526 14716 3834 14736
rect 3526 14714 3532 14716
rect 3588 14714 3612 14716
rect 3668 14714 3692 14716
rect 3748 14714 3772 14716
rect 3828 14714 3834 14716
rect 3588 14662 3590 14714
rect 3770 14662 3772 14714
rect 3526 14660 3532 14662
rect 3588 14660 3612 14662
rect 3668 14660 3692 14662
rect 3748 14660 3772 14662
rect 3828 14660 3834 14662
rect 3526 14640 3834 14660
rect 6102 14172 6410 14192
rect 6102 14170 6108 14172
rect 6164 14170 6188 14172
rect 6244 14170 6268 14172
rect 6324 14170 6348 14172
rect 6404 14170 6410 14172
rect 6164 14118 6166 14170
rect 6346 14118 6348 14170
rect 6102 14116 6108 14118
rect 6164 14116 6188 14118
rect 6244 14116 6268 14118
rect 6324 14116 6348 14118
rect 6404 14116 6410 14118
rect 6102 14096 6410 14116
rect 3526 13628 3834 13648
rect 3526 13626 3532 13628
rect 3588 13626 3612 13628
rect 3668 13626 3692 13628
rect 3748 13626 3772 13628
rect 3828 13626 3834 13628
rect 3588 13574 3590 13626
rect 3770 13574 3772 13626
rect 3526 13572 3532 13574
rect 3588 13572 3612 13574
rect 3668 13572 3692 13574
rect 3748 13572 3772 13574
rect 3828 13572 3834 13574
rect 3526 13552 3834 13572
rect 6102 13084 6410 13104
rect 6102 13082 6108 13084
rect 6164 13082 6188 13084
rect 6244 13082 6268 13084
rect 6324 13082 6348 13084
rect 6404 13082 6410 13084
rect 6164 13030 6166 13082
rect 6346 13030 6348 13082
rect 6102 13028 6108 13030
rect 6164 13028 6188 13030
rect 6244 13028 6268 13030
rect 6324 13028 6348 13030
rect 6404 13028 6410 13030
rect 6102 13008 6410 13028
rect 3526 12540 3834 12560
rect 3526 12538 3532 12540
rect 3588 12538 3612 12540
rect 3668 12538 3692 12540
rect 3748 12538 3772 12540
rect 3828 12538 3834 12540
rect 3588 12486 3590 12538
rect 3770 12486 3772 12538
rect 3526 12484 3532 12486
rect 3588 12484 3612 12486
rect 3668 12484 3692 12486
rect 3748 12484 3772 12486
rect 3828 12484 3834 12486
rect 3526 12464 3834 12484
rect 6102 11996 6410 12016
rect 6102 11994 6108 11996
rect 6164 11994 6188 11996
rect 6244 11994 6268 11996
rect 6324 11994 6348 11996
rect 6404 11994 6410 11996
rect 6164 11942 6166 11994
rect 6346 11942 6348 11994
rect 6102 11940 6108 11942
rect 6164 11940 6188 11942
rect 6244 11940 6268 11942
rect 6324 11940 6348 11942
rect 6404 11940 6410 11942
rect 6102 11920 6410 11940
rect 3526 11452 3834 11472
rect 3526 11450 3532 11452
rect 3588 11450 3612 11452
rect 3668 11450 3692 11452
rect 3748 11450 3772 11452
rect 3828 11450 3834 11452
rect 3588 11398 3590 11450
rect 3770 11398 3772 11450
rect 3526 11396 3532 11398
rect 3588 11396 3612 11398
rect 3668 11396 3692 11398
rect 3748 11396 3772 11398
rect 3828 11396 3834 11398
rect 3526 11376 3834 11396
rect 6102 10908 6410 10928
rect 6102 10906 6108 10908
rect 6164 10906 6188 10908
rect 6244 10906 6268 10908
rect 6324 10906 6348 10908
rect 6404 10906 6410 10908
rect 6164 10854 6166 10906
rect 6346 10854 6348 10906
rect 6102 10852 6108 10854
rect 6164 10852 6188 10854
rect 6244 10852 6268 10854
rect 6324 10852 6348 10854
rect 6404 10852 6410 10854
rect 6102 10832 6410 10852
rect 3526 10364 3834 10384
rect 3526 10362 3532 10364
rect 3588 10362 3612 10364
rect 3668 10362 3692 10364
rect 3748 10362 3772 10364
rect 3828 10362 3834 10364
rect 3588 10310 3590 10362
rect 3770 10310 3772 10362
rect 3526 10308 3532 10310
rect 3588 10308 3612 10310
rect 3668 10308 3692 10310
rect 3748 10308 3772 10310
rect 3828 10308 3834 10310
rect 3526 10288 3834 10308
rect 6102 9820 6410 9840
rect 6102 9818 6108 9820
rect 6164 9818 6188 9820
rect 6244 9818 6268 9820
rect 6324 9818 6348 9820
rect 6404 9818 6410 9820
rect 6164 9766 6166 9818
rect 6346 9766 6348 9818
rect 6102 9764 6108 9766
rect 6164 9764 6188 9766
rect 6244 9764 6268 9766
rect 6324 9764 6348 9766
rect 6404 9764 6410 9766
rect 6102 9744 6410 9764
rect 3526 9276 3834 9296
rect 3526 9274 3532 9276
rect 3588 9274 3612 9276
rect 3668 9274 3692 9276
rect 3748 9274 3772 9276
rect 3828 9274 3834 9276
rect 3588 9222 3590 9274
rect 3770 9222 3772 9274
rect 3526 9220 3532 9222
rect 3588 9220 3612 9222
rect 3668 9220 3692 9222
rect 3748 9220 3772 9222
rect 3828 9220 3834 9222
rect 3526 9200 3834 9220
rect 6102 8732 6410 8752
rect 6102 8730 6108 8732
rect 6164 8730 6188 8732
rect 6244 8730 6268 8732
rect 6324 8730 6348 8732
rect 6404 8730 6410 8732
rect 6164 8678 6166 8730
rect 6346 8678 6348 8730
rect 6102 8676 6108 8678
rect 6164 8676 6188 8678
rect 6244 8676 6268 8678
rect 6324 8676 6348 8678
rect 6404 8676 6410 8678
rect 6102 8656 6410 8676
rect 3526 8188 3834 8208
rect 3526 8186 3532 8188
rect 3588 8186 3612 8188
rect 3668 8186 3692 8188
rect 3748 8186 3772 8188
rect 3828 8186 3834 8188
rect 3588 8134 3590 8186
rect 3770 8134 3772 8186
rect 3526 8132 3532 8134
rect 3588 8132 3612 8134
rect 3668 8132 3692 8134
rect 3748 8132 3772 8134
rect 3828 8132 3834 8134
rect 3526 8112 3834 8132
rect 6102 7644 6410 7664
rect 6102 7642 6108 7644
rect 6164 7642 6188 7644
rect 6244 7642 6268 7644
rect 6324 7642 6348 7644
rect 6404 7642 6410 7644
rect 6164 7590 6166 7642
rect 6346 7590 6348 7642
rect 6102 7588 6108 7590
rect 6164 7588 6188 7590
rect 6244 7588 6268 7590
rect 6324 7588 6348 7590
rect 6404 7588 6410 7590
rect 6102 7568 6410 7588
rect 3526 7100 3834 7120
rect 3526 7098 3532 7100
rect 3588 7098 3612 7100
rect 3668 7098 3692 7100
rect 3748 7098 3772 7100
rect 3828 7098 3834 7100
rect 3588 7046 3590 7098
rect 3770 7046 3772 7098
rect 3526 7044 3532 7046
rect 3588 7044 3612 7046
rect 3668 7044 3692 7046
rect 3748 7044 3772 7046
rect 3828 7044 3834 7046
rect 3526 7024 3834 7044
rect 7760 6914 7788 17002
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7668 6886 7788 6914
rect 6102 6556 6410 6576
rect 6102 6554 6108 6556
rect 6164 6554 6188 6556
rect 6244 6554 6268 6556
rect 6324 6554 6348 6556
rect 6404 6554 6410 6556
rect 6164 6502 6166 6554
rect 6346 6502 6348 6554
rect 6102 6500 6108 6502
rect 6164 6500 6188 6502
rect 6244 6500 6268 6502
rect 6324 6500 6348 6502
rect 6404 6500 6410 6502
rect 6102 6480 6410 6500
rect 3526 6012 3834 6032
rect 3526 6010 3532 6012
rect 3588 6010 3612 6012
rect 3668 6010 3692 6012
rect 3748 6010 3772 6012
rect 3828 6010 3834 6012
rect 3588 5958 3590 6010
rect 3770 5958 3772 6010
rect 3526 5956 3532 5958
rect 3588 5956 3612 5958
rect 3668 5956 3692 5958
rect 3748 5956 3772 5958
rect 3828 5956 3834 5958
rect 3526 5936 3834 5956
rect 6102 5468 6410 5488
rect 6102 5466 6108 5468
rect 6164 5466 6188 5468
rect 6244 5466 6268 5468
rect 6324 5466 6348 5468
rect 6404 5466 6410 5468
rect 6164 5414 6166 5466
rect 6346 5414 6348 5466
rect 6102 5412 6108 5414
rect 6164 5412 6188 5414
rect 6244 5412 6268 5414
rect 6324 5412 6348 5414
rect 6404 5412 6410 5414
rect 6102 5392 6410 5412
rect 7668 5234 7696 6886
rect 7852 5234 7880 16934
rect 8678 16892 8986 16912
rect 8678 16890 8684 16892
rect 8740 16890 8764 16892
rect 8820 16890 8844 16892
rect 8900 16890 8924 16892
rect 8980 16890 8986 16892
rect 8740 16838 8742 16890
rect 8922 16838 8924 16890
rect 8678 16836 8684 16838
rect 8740 16836 8764 16838
rect 8820 16836 8844 16838
rect 8900 16836 8924 16838
rect 8980 16836 8986 16838
rect 8678 16816 8986 16836
rect 13830 16892 14138 16912
rect 13830 16890 13836 16892
rect 13892 16890 13916 16892
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14138 16892
rect 13892 16838 13894 16890
rect 14074 16838 14076 16890
rect 13830 16836 13836 16838
rect 13892 16836 13916 16838
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14138 16838
rect 13830 16816 14138 16836
rect 11254 16348 11562 16368
rect 11254 16346 11260 16348
rect 11316 16346 11340 16348
rect 11396 16346 11420 16348
rect 11476 16346 11500 16348
rect 11556 16346 11562 16348
rect 11316 16294 11318 16346
rect 11498 16294 11500 16346
rect 11254 16292 11260 16294
rect 11316 16292 11340 16294
rect 11396 16292 11420 16294
rect 11476 16292 11500 16294
rect 11556 16292 11562 16294
rect 11254 16272 11562 16292
rect 8678 15804 8986 15824
rect 8678 15802 8684 15804
rect 8740 15802 8764 15804
rect 8820 15802 8844 15804
rect 8900 15802 8924 15804
rect 8980 15802 8986 15804
rect 8740 15750 8742 15802
rect 8922 15750 8924 15802
rect 8678 15748 8684 15750
rect 8740 15748 8764 15750
rect 8820 15748 8844 15750
rect 8900 15748 8924 15750
rect 8980 15748 8986 15750
rect 8678 15728 8986 15748
rect 13830 15804 14138 15824
rect 13830 15802 13836 15804
rect 13892 15802 13916 15804
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14138 15804
rect 13892 15750 13894 15802
rect 14074 15750 14076 15802
rect 13830 15748 13836 15750
rect 13892 15748 13916 15750
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14138 15750
rect 13830 15728 14138 15748
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8678 14716 8986 14736
rect 8678 14714 8684 14716
rect 8740 14714 8764 14716
rect 8820 14714 8844 14716
rect 8900 14714 8924 14716
rect 8980 14714 8986 14716
rect 8740 14662 8742 14714
rect 8922 14662 8924 14714
rect 8678 14660 8684 14662
rect 8740 14660 8764 14662
rect 8820 14660 8844 14662
rect 8900 14660 8924 14662
rect 8980 14660 8986 14662
rect 8678 14640 8986 14660
rect 8678 13628 8986 13648
rect 8678 13626 8684 13628
rect 8740 13626 8764 13628
rect 8820 13626 8844 13628
rect 8900 13626 8924 13628
rect 8980 13626 8986 13628
rect 8740 13574 8742 13626
rect 8922 13574 8924 13626
rect 8678 13572 8684 13574
rect 8740 13572 8764 13574
rect 8820 13572 8844 13574
rect 8900 13572 8924 13574
rect 8980 13572 8986 13574
rect 8678 13552 8986 13572
rect 8678 12540 8986 12560
rect 8678 12538 8684 12540
rect 8740 12538 8764 12540
rect 8820 12538 8844 12540
rect 8900 12538 8924 12540
rect 8980 12538 8986 12540
rect 8740 12486 8742 12538
rect 8922 12486 8924 12538
rect 8678 12484 8684 12486
rect 8740 12484 8764 12486
rect 8820 12484 8844 12486
rect 8900 12484 8924 12486
rect 8980 12484 8986 12486
rect 8678 12464 8986 12484
rect 8678 11452 8986 11472
rect 8678 11450 8684 11452
rect 8740 11450 8764 11452
rect 8820 11450 8844 11452
rect 8900 11450 8924 11452
rect 8980 11450 8986 11452
rect 8740 11398 8742 11450
rect 8922 11398 8924 11450
rect 8678 11396 8684 11398
rect 8740 11396 8764 11398
rect 8820 11396 8844 11398
rect 8900 11396 8924 11398
rect 8980 11396 8986 11398
rect 8678 11376 8986 11396
rect 8678 10364 8986 10384
rect 8678 10362 8684 10364
rect 8740 10362 8764 10364
rect 8820 10362 8844 10364
rect 8900 10362 8924 10364
rect 8980 10362 8986 10364
rect 8740 10310 8742 10362
rect 8922 10310 8924 10362
rect 8678 10308 8684 10310
rect 8740 10308 8764 10310
rect 8820 10308 8844 10310
rect 8900 10308 8924 10310
rect 8980 10308 8986 10310
rect 8678 10288 8986 10308
rect 8678 9276 8986 9296
rect 8678 9274 8684 9276
rect 8740 9274 8764 9276
rect 8820 9274 8844 9276
rect 8900 9274 8924 9276
rect 8980 9274 8986 9276
rect 8740 9222 8742 9274
rect 8922 9222 8924 9274
rect 8678 9220 8684 9222
rect 8740 9220 8764 9222
rect 8820 9220 8844 9222
rect 8900 9220 8924 9222
rect 8980 9220 8986 9222
rect 8678 9200 8986 9220
rect 8678 8188 8986 8208
rect 8678 8186 8684 8188
rect 8740 8186 8764 8188
rect 8820 8186 8844 8188
rect 8900 8186 8924 8188
rect 8980 8186 8986 8188
rect 8740 8134 8742 8186
rect 8922 8134 8924 8186
rect 8678 8132 8684 8134
rect 8740 8132 8764 8134
rect 8820 8132 8844 8134
rect 8900 8132 8924 8134
rect 8980 8132 8986 8134
rect 8678 8112 8986 8132
rect 8678 7100 8986 7120
rect 8678 7098 8684 7100
rect 8740 7098 8764 7100
rect 8820 7098 8844 7100
rect 8900 7098 8924 7100
rect 8980 7098 8986 7100
rect 8740 7046 8742 7098
rect 8922 7046 8924 7098
rect 8678 7044 8684 7046
rect 8740 7044 8764 7046
rect 8820 7044 8844 7046
rect 8900 7044 8924 7046
rect 8980 7044 8986 7046
rect 8678 7024 8986 7044
rect 8678 6012 8986 6032
rect 8678 6010 8684 6012
rect 8740 6010 8764 6012
rect 8820 6010 8844 6012
rect 8900 6010 8924 6012
rect 8980 6010 8986 6012
rect 8740 5958 8742 6010
rect 8922 5958 8924 6010
rect 8678 5956 8684 5958
rect 8740 5956 8764 5958
rect 8820 5956 8844 5958
rect 8900 5956 8924 5958
rect 8980 5956 8986 5958
rect 8678 5936 8986 5956
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 3526 4924 3834 4944
rect 3526 4922 3532 4924
rect 3588 4922 3612 4924
rect 3668 4922 3692 4924
rect 3748 4922 3772 4924
rect 3828 4922 3834 4924
rect 3588 4870 3590 4922
rect 3770 4870 3772 4922
rect 3526 4868 3532 4870
rect 3588 4868 3612 4870
rect 3668 4868 3692 4870
rect 3748 4868 3772 4870
rect 3828 4868 3834 4870
rect 3526 4848 3834 4868
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6102 4380 6410 4400
rect 6102 4378 6108 4380
rect 6164 4378 6188 4380
rect 6244 4378 6268 4380
rect 6324 4378 6348 4380
rect 6404 4378 6410 4380
rect 6164 4326 6166 4378
rect 6346 4326 6348 4378
rect 6102 4324 6108 4326
rect 6164 4324 6188 4326
rect 6244 4324 6268 4326
rect 6324 4324 6348 4326
rect 6404 4324 6410 4326
rect 6102 4304 6410 4324
rect 6472 4162 6500 4558
rect 6840 4486 6868 5034
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4690 6960 4966
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6380 4134 6500 4162
rect 6380 4078 6408 4134
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 3526 3836 3834 3856
rect 3526 3834 3532 3836
rect 3588 3834 3612 3836
rect 3668 3834 3692 3836
rect 3748 3834 3772 3836
rect 3828 3834 3834 3836
rect 3588 3782 3590 3834
rect 3770 3782 3772 3834
rect 3526 3780 3532 3782
rect 3588 3780 3612 3782
rect 3668 3780 3692 3782
rect 3748 3780 3772 3782
rect 3828 3780 3834 3782
rect 3526 3760 3834 3780
rect 6380 3534 6408 4014
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 5552 3398 5580 3470
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5920 3194 5948 3470
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5920 2854 5948 3130
rect 6012 3126 6040 3470
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6102 3292 6410 3312
rect 6102 3290 6108 3292
rect 6164 3290 6188 3292
rect 6244 3290 6268 3292
rect 6324 3290 6348 3292
rect 6404 3290 6410 3292
rect 6164 3238 6166 3290
rect 6346 3238 6348 3290
rect 6102 3236 6108 3238
rect 6164 3236 6188 3238
rect 6244 3236 6268 3238
rect 6324 3236 6348 3238
rect 6404 3236 6410 3238
rect 6102 3216 6410 3236
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 3526 2748 3834 2768
rect 3526 2746 3532 2748
rect 3588 2746 3612 2748
rect 3668 2746 3692 2748
rect 3748 2746 3772 2748
rect 3828 2746 3834 2748
rect 3588 2694 3590 2746
rect 3770 2694 3772 2746
rect 3526 2692 3532 2694
rect 3588 2692 3612 2694
rect 3668 2692 3692 2694
rect 3748 2692 3772 2694
rect 3828 2692 3834 2694
rect 3526 2672 3834 2692
rect 6564 2446 6592 3334
rect 6656 2650 6684 4014
rect 6748 3058 6776 4014
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6840 2582 6868 4422
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6932 2394 6960 2790
rect 7024 2514 7052 3674
rect 7668 3398 7696 5170
rect 8220 4622 8248 5170
rect 8678 4924 8986 4944
rect 8678 4922 8684 4924
rect 8740 4922 8764 4924
rect 8820 4922 8844 4924
rect 8900 4922 8924 4924
rect 8980 4922 8986 4924
rect 8740 4870 8742 4922
rect 8922 4870 8924 4922
rect 8678 4868 8684 4870
rect 8740 4868 8764 4870
rect 8820 4868 8844 4870
rect 8900 4868 8924 4870
rect 8980 4868 8986 4870
rect 8678 4848 8986 4868
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8036 4214 8064 4558
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7944 3398 7972 3538
rect 8036 3466 8064 4150
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3738 8156 3878
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7300 2650 7328 2926
rect 7944 2774 7972 3334
rect 8036 3126 8064 3402
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7852 2746 7972 2774
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7852 2446 7880 2746
rect 8220 2446 8248 4558
rect 9048 4214 9076 15302
rect 11254 15260 11562 15280
rect 11254 15258 11260 15260
rect 11316 15258 11340 15260
rect 11396 15258 11420 15260
rect 11476 15258 11500 15260
rect 11556 15258 11562 15260
rect 11316 15206 11318 15258
rect 11498 15206 11500 15258
rect 11254 15204 11260 15206
rect 11316 15204 11340 15206
rect 11396 15204 11420 15206
rect 11476 15204 11500 15206
rect 11556 15204 11562 15206
rect 11254 15184 11562 15204
rect 13830 14716 14138 14736
rect 13830 14714 13836 14716
rect 13892 14714 13916 14716
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14138 14716
rect 13892 14662 13894 14714
rect 14074 14662 14076 14714
rect 13830 14660 13836 14662
rect 13892 14660 13916 14662
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14138 14662
rect 13830 14640 14138 14660
rect 11254 14172 11562 14192
rect 11254 14170 11260 14172
rect 11316 14170 11340 14172
rect 11396 14170 11420 14172
rect 11476 14170 11500 14172
rect 11556 14170 11562 14172
rect 11316 14118 11318 14170
rect 11498 14118 11500 14170
rect 11254 14116 11260 14118
rect 11316 14116 11340 14118
rect 11396 14116 11420 14118
rect 11476 14116 11500 14118
rect 11556 14116 11562 14118
rect 11254 14096 11562 14116
rect 13830 13628 14138 13648
rect 13830 13626 13836 13628
rect 13892 13626 13916 13628
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14138 13628
rect 13892 13574 13894 13626
rect 14074 13574 14076 13626
rect 13830 13572 13836 13574
rect 13892 13572 13916 13574
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14138 13574
rect 13830 13552 14138 13572
rect 11254 13084 11562 13104
rect 11254 13082 11260 13084
rect 11316 13082 11340 13084
rect 11396 13082 11420 13084
rect 11476 13082 11500 13084
rect 11556 13082 11562 13084
rect 11316 13030 11318 13082
rect 11498 13030 11500 13082
rect 11254 13028 11260 13030
rect 11316 13028 11340 13030
rect 11396 13028 11420 13030
rect 11476 13028 11500 13030
rect 11556 13028 11562 13030
rect 11254 13008 11562 13028
rect 13830 12540 14138 12560
rect 13830 12538 13836 12540
rect 13892 12538 13916 12540
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14138 12540
rect 13892 12486 13894 12538
rect 14074 12486 14076 12538
rect 13830 12484 13836 12486
rect 13892 12484 13916 12486
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14138 12486
rect 13830 12464 14138 12484
rect 11254 11996 11562 12016
rect 11254 11994 11260 11996
rect 11316 11994 11340 11996
rect 11396 11994 11420 11996
rect 11476 11994 11500 11996
rect 11556 11994 11562 11996
rect 11316 11942 11318 11994
rect 11498 11942 11500 11994
rect 11254 11940 11260 11942
rect 11316 11940 11340 11942
rect 11396 11940 11420 11942
rect 11476 11940 11500 11942
rect 11556 11940 11562 11942
rect 11254 11920 11562 11940
rect 13830 11452 14138 11472
rect 13830 11450 13836 11452
rect 13892 11450 13916 11452
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14138 11452
rect 13892 11398 13894 11450
rect 14074 11398 14076 11450
rect 13830 11396 13836 11398
rect 13892 11396 13916 11398
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14138 11398
rect 13830 11376 14138 11396
rect 11254 10908 11562 10928
rect 11254 10906 11260 10908
rect 11316 10906 11340 10908
rect 11396 10906 11420 10908
rect 11476 10906 11500 10908
rect 11556 10906 11562 10908
rect 11316 10854 11318 10906
rect 11498 10854 11500 10906
rect 11254 10852 11260 10854
rect 11316 10852 11340 10854
rect 11396 10852 11420 10854
rect 11476 10852 11500 10854
rect 11556 10852 11562 10854
rect 11254 10832 11562 10852
rect 13830 10364 14138 10384
rect 13830 10362 13836 10364
rect 13892 10362 13916 10364
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14138 10364
rect 13892 10310 13894 10362
rect 14074 10310 14076 10362
rect 13830 10308 13836 10310
rect 13892 10308 13916 10310
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14138 10310
rect 13830 10288 14138 10308
rect 11254 9820 11562 9840
rect 11254 9818 11260 9820
rect 11316 9818 11340 9820
rect 11396 9818 11420 9820
rect 11476 9818 11500 9820
rect 11556 9818 11562 9820
rect 11316 9766 11318 9818
rect 11498 9766 11500 9818
rect 11254 9764 11260 9766
rect 11316 9764 11340 9766
rect 11396 9764 11420 9766
rect 11476 9764 11500 9766
rect 11556 9764 11562 9766
rect 11254 9744 11562 9764
rect 13830 9276 14138 9296
rect 13830 9274 13836 9276
rect 13892 9274 13916 9276
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14138 9276
rect 13892 9222 13894 9274
rect 14074 9222 14076 9274
rect 13830 9220 13836 9222
rect 13892 9220 13916 9222
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14138 9222
rect 13830 9200 14138 9220
rect 11254 8732 11562 8752
rect 11254 8730 11260 8732
rect 11316 8730 11340 8732
rect 11396 8730 11420 8732
rect 11476 8730 11500 8732
rect 11556 8730 11562 8732
rect 11316 8678 11318 8730
rect 11498 8678 11500 8730
rect 11254 8676 11260 8678
rect 11316 8676 11340 8678
rect 11396 8676 11420 8678
rect 11476 8676 11500 8678
rect 11556 8676 11562 8678
rect 11254 8656 11562 8676
rect 13830 8188 14138 8208
rect 13830 8186 13836 8188
rect 13892 8186 13916 8188
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14138 8188
rect 13892 8134 13894 8186
rect 14074 8134 14076 8186
rect 13830 8132 13836 8134
rect 13892 8132 13916 8134
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14138 8134
rect 13830 8112 14138 8132
rect 11254 7644 11562 7664
rect 11254 7642 11260 7644
rect 11316 7642 11340 7644
rect 11396 7642 11420 7644
rect 11476 7642 11500 7644
rect 11556 7642 11562 7644
rect 11316 7590 11318 7642
rect 11498 7590 11500 7642
rect 11254 7588 11260 7590
rect 11316 7588 11340 7590
rect 11396 7588 11420 7590
rect 11476 7588 11500 7590
rect 11556 7588 11562 7590
rect 11254 7568 11562 7588
rect 13830 7100 14138 7120
rect 13830 7098 13836 7100
rect 13892 7098 13916 7100
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14138 7100
rect 13892 7046 13894 7098
rect 14074 7046 14076 7098
rect 13830 7044 13836 7046
rect 13892 7044 13916 7046
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14138 7046
rect 13830 7024 14138 7044
rect 11254 6556 11562 6576
rect 11254 6554 11260 6556
rect 11316 6554 11340 6556
rect 11396 6554 11420 6556
rect 11476 6554 11500 6556
rect 11556 6554 11562 6556
rect 11316 6502 11318 6554
rect 11498 6502 11500 6554
rect 11254 6500 11260 6502
rect 11316 6500 11340 6502
rect 11396 6500 11420 6502
rect 11476 6500 11500 6502
rect 11556 6500 11562 6502
rect 11254 6480 11562 6500
rect 13830 6012 14138 6032
rect 13830 6010 13836 6012
rect 13892 6010 13916 6012
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14138 6012
rect 13892 5958 13894 6010
rect 14074 5958 14076 6010
rect 13830 5956 13836 5958
rect 13892 5956 13916 5958
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14138 5958
rect 13830 5936 14138 5956
rect 11254 5468 11562 5488
rect 11254 5466 11260 5468
rect 11316 5466 11340 5468
rect 11396 5466 11420 5468
rect 11476 5466 11500 5468
rect 11556 5466 11562 5468
rect 11316 5414 11318 5466
rect 11498 5414 11500 5466
rect 11254 5412 11260 5414
rect 11316 5412 11340 5414
rect 11396 5412 11420 5414
rect 11476 5412 11500 5414
rect 11556 5412 11562 5414
rect 11254 5392 11562 5412
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8678 3836 8986 3856
rect 8678 3834 8684 3836
rect 8740 3834 8764 3836
rect 8820 3834 8844 3836
rect 8900 3834 8924 3836
rect 8980 3834 8986 3836
rect 8740 3782 8742 3834
rect 8922 3782 8924 3834
rect 8678 3780 8684 3782
rect 8740 3780 8764 3782
rect 8820 3780 8844 3782
rect 8900 3780 8924 3782
rect 8980 3780 8986 3782
rect 8678 3760 8986 3780
rect 9140 3738 9168 4626
rect 9324 4622 9352 4966
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9232 3194 9260 4558
rect 9324 4214 9352 4558
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 8678 2748 8986 2768
rect 8678 2746 8684 2748
rect 8740 2746 8764 2748
rect 8820 2746 8844 2748
rect 8900 2746 8924 2748
rect 8980 2746 8986 2748
rect 8740 2694 8742 2746
rect 8922 2694 8924 2746
rect 8678 2692 8684 2694
rect 8740 2692 8764 2694
rect 8820 2692 8844 2694
rect 8900 2692 8924 2694
rect 8980 2692 8986 2694
rect 8678 2672 8986 2692
rect 9232 2514 9260 3130
rect 9324 2582 9352 4150
rect 9692 4078 9720 4966
rect 13830 4924 14138 4944
rect 13830 4922 13836 4924
rect 13892 4922 13916 4924
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14138 4924
rect 13892 4870 13894 4922
rect 14074 4870 14076 4922
rect 13830 4868 13836 4870
rect 13892 4868 13916 4870
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14138 4870
rect 13830 4848 14138 4868
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 12164 4548 12216 4554
rect 12164 4490 12216 4496
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3058 10364 3878
rect 10428 3602 10456 4422
rect 10704 3602 10732 4422
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10704 3194 10732 3538
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10796 2582 10824 4490
rect 11254 4380 11562 4400
rect 11254 4378 11260 4380
rect 11316 4378 11340 4380
rect 11396 4378 11420 4380
rect 11476 4378 11500 4380
rect 11556 4378 11562 4380
rect 11316 4326 11318 4378
rect 11498 4326 11500 4378
rect 11254 4324 11260 4326
rect 11316 4324 11340 4326
rect 11396 4324 11420 4326
rect 11476 4324 11500 4326
rect 11556 4324 11562 4326
rect 11254 4304 11562 4324
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 2650 10916 4014
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3602 11468 3878
rect 11808 3738 11836 4082
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11254 3292 11562 3312
rect 11254 3290 11260 3292
rect 11316 3290 11340 3292
rect 11396 3290 11420 3292
rect 11476 3290 11500 3292
rect 11556 3290 11562 3292
rect 11316 3238 11318 3290
rect 11498 3238 11500 3290
rect 11254 3236 11260 3238
rect 11316 3236 11340 3238
rect 11396 3236 11420 3238
rect 11476 3236 11500 3238
rect 11556 3236 11562 3238
rect 11254 3216 11562 3236
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 11808 2446 11836 3674
rect 12084 3126 12112 3878
rect 12176 3466 12204 4490
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 4146 12388 4422
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12176 3194 12204 3402
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 12360 2582 12388 4082
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12452 3398 12480 4014
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12452 2446 12480 3334
rect 13004 2854 13032 3878
rect 13830 3836 14138 3856
rect 13830 3834 13836 3836
rect 13892 3834 13916 3836
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14138 3836
rect 13892 3782 13894 3834
rect 14074 3782 14076 3834
rect 13830 3780 13836 3782
rect 13892 3780 13916 3782
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14138 3782
rect 13830 3760 14138 3780
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 13830 2748 14138 2768
rect 13830 2746 13836 2748
rect 13892 2746 13916 2748
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14138 2748
rect 13892 2694 13894 2746
rect 14074 2694 14076 2746
rect 13830 2692 13836 2694
rect 13892 2692 13916 2694
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14138 2694
rect 13830 2672 14138 2692
rect 15672 2446 15700 2790
rect 7104 2440 7156 2446
rect 6932 2388 7104 2394
rect 7840 2440 7892 2446
rect 6932 2382 7156 2388
rect 7668 2400 7840 2428
rect 1124 2372 1176 2378
rect 1124 2314 1176 2320
rect 3332 2372 3384 2378
rect 3332 2314 3384 2320
rect 5540 2372 5592 2378
rect 6932 2366 7144 2382
rect 5540 2314 5592 2320
rect 1136 800 1164 2314
rect 3344 800 3372 2314
rect 5552 800 5580 2314
rect 7668 2310 7696 2400
rect 7840 2382 7892 2388
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 10784 2372 10836 2378
rect 10784 2314 10836 2320
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 6102 2204 6410 2224
rect 6102 2202 6108 2204
rect 6164 2202 6188 2204
rect 6244 2202 6268 2204
rect 6324 2202 6348 2204
rect 6404 2202 6410 2204
rect 6164 2150 6166 2202
rect 6346 2150 6348 2202
rect 6102 2148 6108 2150
rect 6164 2148 6188 2150
rect 6244 2148 6268 2150
rect 6324 2148 6348 2150
rect 6404 2148 6410 2150
rect 6102 2128 6410 2148
rect 7760 800 7788 2246
rect 10796 898 10824 2314
rect 11254 2204 11562 2224
rect 11254 2202 11260 2204
rect 11316 2202 11340 2204
rect 11396 2202 11420 2204
rect 11476 2202 11500 2204
rect 11556 2202 11562 2204
rect 11316 2150 11318 2202
rect 11498 2150 11500 2202
rect 11254 2148 11260 2150
rect 11316 2148 11340 2150
rect 11396 2148 11420 2150
rect 11476 2148 11500 2150
rect 11556 2148 11562 2150
rect 11254 2128 11562 2148
rect 9968 870 10088 898
rect 9968 800 9996 870
rect 1122 0 1178 800
rect 3330 0 3386 800
rect 5538 0 5594 800
rect 7746 0 7802 800
rect 9954 0 10010 800
rect 10060 762 10088 870
rect 10336 870 10824 898
rect 10336 762 10364 870
rect 12176 800 12204 2314
rect 12452 2310 12480 2382
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 14384 800 14412 2314
rect 16592 800 16620 2314
rect 10060 734 10364 762
rect 12162 0 12218 800
rect 14370 0 14426 800
rect 16578 0 16634 800
<< via2 >>
rect 6108 17434 6164 17436
rect 6188 17434 6244 17436
rect 6268 17434 6324 17436
rect 6348 17434 6404 17436
rect 6108 17382 6154 17434
rect 6154 17382 6164 17434
rect 6188 17382 6218 17434
rect 6218 17382 6230 17434
rect 6230 17382 6244 17434
rect 6268 17382 6282 17434
rect 6282 17382 6294 17434
rect 6294 17382 6324 17434
rect 6348 17382 6358 17434
rect 6358 17382 6404 17434
rect 6108 17380 6164 17382
rect 6188 17380 6244 17382
rect 6268 17380 6324 17382
rect 6348 17380 6404 17382
rect 3532 16890 3588 16892
rect 3612 16890 3668 16892
rect 3692 16890 3748 16892
rect 3772 16890 3828 16892
rect 3532 16838 3578 16890
rect 3578 16838 3588 16890
rect 3612 16838 3642 16890
rect 3642 16838 3654 16890
rect 3654 16838 3668 16890
rect 3692 16838 3706 16890
rect 3706 16838 3718 16890
rect 3718 16838 3748 16890
rect 3772 16838 3782 16890
rect 3782 16838 3828 16890
rect 3532 16836 3588 16838
rect 3612 16836 3668 16838
rect 3692 16836 3748 16838
rect 3772 16836 3828 16838
rect 6108 16346 6164 16348
rect 6188 16346 6244 16348
rect 6268 16346 6324 16348
rect 6348 16346 6404 16348
rect 6108 16294 6154 16346
rect 6154 16294 6164 16346
rect 6188 16294 6218 16346
rect 6218 16294 6230 16346
rect 6230 16294 6244 16346
rect 6268 16294 6282 16346
rect 6282 16294 6294 16346
rect 6294 16294 6324 16346
rect 6348 16294 6358 16346
rect 6358 16294 6404 16346
rect 6108 16292 6164 16294
rect 6188 16292 6244 16294
rect 6268 16292 6324 16294
rect 6348 16292 6404 16294
rect 3532 15802 3588 15804
rect 3612 15802 3668 15804
rect 3692 15802 3748 15804
rect 3772 15802 3828 15804
rect 3532 15750 3578 15802
rect 3578 15750 3588 15802
rect 3612 15750 3642 15802
rect 3642 15750 3654 15802
rect 3654 15750 3668 15802
rect 3692 15750 3706 15802
rect 3706 15750 3718 15802
rect 3718 15750 3748 15802
rect 3772 15750 3782 15802
rect 3782 15750 3828 15802
rect 3532 15748 3588 15750
rect 3612 15748 3668 15750
rect 3692 15748 3748 15750
rect 3772 15748 3828 15750
rect 11260 17434 11316 17436
rect 11340 17434 11396 17436
rect 11420 17434 11476 17436
rect 11500 17434 11556 17436
rect 11260 17382 11306 17434
rect 11306 17382 11316 17434
rect 11340 17382 11370 17434
rect 11370 17382 11382 17434
rect 11382 17382 11396 17434
rect 11420 17382 11434 17434
rect 11434 17382 11446 17434
rect 11446 17382 11476 17434
rect 11500 17382 11510 17434
rect 11510 17382 11556 17434
rect 11260 17380 11316 17382
rect 11340 17380 11396 17382
rect 11420 17380 11476 17382
rect 11500 17380 11556 17382
rect 6108 15258 6164 15260
rect 6188 15258 6244 15260
rect 6268 15258 6324 15260
rect 6348 15258 6404 15260
rect 6108 15206 6154 15258
rect 6154 15206 6164 15258
rect 6188 15206 6218 15258
rect 6218 15206 6230 15258
rect 6230 15206 6244 15258
rect 6268 15206 6282 15258
rect 6282 15206 6294 15258
rect 6294 15206 6324 15258
rect 6348 15206 6358 15258
rect 6358 15206 6404 15258
rect 6108 15204 6164 15206
rect 6188 15204 6244 15206
rect 6268 15204 6324 15206
rect 6348 15204 6404 15206
rect 3532 14714 3588 14716
rect 3612 14714 3668 14716
rect 3692 14714 3748 14716
rect 3772 14714 3828 14716
rect 3532 14662 3578 14714
rect 3578 14662 3588 14714
rect 3612 14662 3642 14714
rect 3642 14662 3654 14714
rect 3654 14662 3668 14714
rect 3692 14662 3706 14714
rect 3706 14662 3718 14714
rect 3718 14662 3748 14714
rect 3772 14662 3782 14714
rect 3782 14662 3828 14714
rect 3532 14660 3588 14662
rect 3612 14660 3668 14662
rect 3692 14660 3748 14662
rect 3772 14660 3828 14662
rect 6108 14170 6164 14172
rect 6188 14170 6244 14172
rect 6268 14170 6324 14172
rect 6348 14170 6404 14172
rect 6108 14118 6154 14170
rect 6154 14118 6164 14170
rect 6188 14118 6218 14170
rect 6218 14118 6230 14170
rect 6230 14118 6244 14170
rect 6268 14118 6282 14170
rect 6282 14118 6294 14170
rect 6294 14118 6324 14170
rect 6348 14118 6358 14170
rect 6358 14118 6404 14170
rect 6108 14116 6164 14118
rect 6188 14116 6244 14118
rect 6268 14116 6324 14118
rect 6348 14116 6404 14118
rect 3532 13626 3588 13628
rect 3612 13626 3668 13628
rect 3692 13626 3748 13628
rect 3772 13626 3828 13628
rect 3532 13574 3578 13626
rect 3578 13574 3588 13626
rect 3612 13574 3642 13626
rect 3642 13574 3654 13626
rect 3654 13574 3668 13626
rect 3692 13574 3706 13626
rect 3706 13574 3718 13626
rect 3718 13574 3748 13626
rect 3772 13574 3782 13626
rect 3782 13574 3828 13626
rect 3532 13572 3588 13574
rect 3612 13572 3668 13574
rect 3692 13572 3748 13574
rect 3772 13572 3828 13574
rect 6108 13082 6164 13084
rect 6188 13082 6244 13084
rect 6268 13082 6324 13084
rect 6348 13082 6404 13084
rect 6108 13030 6154 13082
rect 6154 13030 6164 13082
rect 6188 13030 6218 13082
rect 6218 13030 6230 13082
rect 6230 13030 6244 13082
rect 6268 13030 6282 13082
rect 6282 13030 6294 13082
rect 6294 13030 6324 13082
rect 6348 13030 6358 13082
rect 6358 13030 6404 13082
rect 6108 13028 6164 13030
rect 6188 13028 6244 13030
rect 6268 13028 6324 13030
rect 6348 13028 6404 13030
rect 3532 12538 3588 12540
rect 3612 12538 3668 12540
rect 3692 12538 3748 12540
rect 3772 12538 3828 12540
rect 3532 12486 3578 12538
rect 3578 12486 3588 12538
rect 3612 12486 3642 12538
rect 3642 12486 3654 12538
rect 3654 12486 3668 12538
rect 3692 12486 3706 12538
rect 3706 12486 3718 12538
rect 3718 12486 3748 12538
rect 3772 12486 3782 12538
rect 3782 12486 3828 12538
rect 3532 12484 3588 12486
rect 3612 12484 3668 12486
rect 3692 12484 3748 12486
rect 3772 12484 3828 12486
rect 6108 11994 6164 11996
rect 6188 11994 6244 11996
rect 6268 11994 6324 11996
rect 6348 11994 6404 11996
rect 6108 11942 6154 11994
rect 6154 11942 6164 11994
rect 6188 11942 6218 11994
rect 6218 11942 6230 11994
rect 6230 11942 6244 11994
rect 6268 11942 6282 11994
rect 6282 11942 6294 11994
rect 6294 11942 6324 11994
rect 6348 11942 6358 11994
rect 6358 11942 6404 11994
rect 6108 11940 6164 11942
rect 6188 11940 6244 11942
rect 6268 11940 6324 11942
rect 6348 11940 6404 11942
rect 3532 11450 3588 11452
rect 3612 11450 3668 11452
rect 3692 11450 3748 11452
rect 3772 11450 3828 11452
rect 3532 11398 3578 11450
rect 3578 11398 3588 11450
rect 3612 11398 3642 11450
rect 3642 11398 3654 11450
rect 3654 11398 3668 11450
rect 3692 11398 3706 11450
rect 3706 11398 3718 11450
rect 3718 11398 3748 11450
rect 3772 11398 3782 11450
rect 3782 11398 3828 11450
rect 3532 11396 3588 11398
rect 3612 11396 3668 11398
rect 3692 11396 3748 11398
rect 3772 11396 3828 11398
rect 6108 10906 6164 10908
rect 6188 10906 6244 10908
rect 6268 10906 6324 10908
rect 6348 10906 6404 10908
rect 6108 10854 6154 10906
rect 6154 10854 6164 10906
rect 6188 10854 6218 10906
rect 6218 10854 6230 10906
rect 6230 10854 6244 10906
rect 6268 10854 6282 10906
rect 6282 10854 6294 10906
rect 6294 10854 6324 10906
rect 6348 10854 6358 10906
rect 6358 10854 6404 10906
rect 6108 10852 6164 10854
rect 6188 10852 6244 10854
rect 6268 10852 6324 10854
rect 6348 10852 6404 10854
rect 3532 10362 3588 10364
rect 3612 10362 3668 10364
rect 3692 10362 3748 10364
rect 3772 10362 3828 10364
rect 3532 10310 3578 10362
rect 3578 10310 3588 10362
rect 3612 10310 3642 10362
rect 3642 10310 3654 10362
rect 3654 10310 3668 10362
rect 3692 10310 3706 10362
rect 3706 10310 3718 10362
rect 3718 10310 3748 10362
rect 3772 10310 3782 10362
rect 3782 10310 3828 10362
rect 3532 10308 3588 10310
rect 3612 10308 3668 10310
rect 3692 10308 3748 10310
rect 3772 10308 3828 10310
rect 6108 9818 6164 9820
rect 6188 9818 6244 9820
rect 6268 9818 6324 9820
rect 6348 9818 6404 9820
rect 6108 9766 6154 9818
rect 6154 9766 6164 9818
rect 6188 9766 6218 9818
rect 6218 9766 6230 9818
rect 6230 9766 6244 9818
rect 6268 9766 6282 9818
rect 6282 9766 6294 9818
rect 6294 9766 6324 9818
rect 6348 9766 6358 9818
rect 6358 9766 6404 9818
rect 6108 9764 6164 9766
rect 6188 9764 6244 9766
rect 6268 9764 6324 9766
rect 6348 9764 6404 9766
rect 3532 9274 3588 9276
rect 3612 9274 3668 9276
rect 3692 9274 3748 9276
rect 3772 9274 3828 9276
rect 3532 9222 3578 9274
rect 3578 9222 3588 9274
rect 3612 9222 3642 9274
rect 3642 9222 3654 9274
rect 3654 9222 3668 9274
rect 3692 9222 3706 9274
rect 3706 9222 3718 9274
rect 3718 9222 3748 9274
rect 3772 9222 3782 9274
rect 3782 9222 3828 9274
rect 3532 9220 3588 9222
rect 3612 9220 3668 9222
rect 3692 9220 3748 9222
rect 3772 9220 3828 9222
rect 6108 8730 6164 8732
rect 6188 8730 6244 8732
rect 6268 8730 6324 8732
rect 6348 8730 6404 8732
rect 6108 8678 6154 8730
rect 6154 8678 6164 8730
rect 6188 8678 6218 8730
rect 6218 8678 6230 8730
rect 6230 8678 6244 8730
rect 6268 8678 6282 8730
rect 6282 8678 6294 8730
rect 6294 8678 6324 8730
rect 6348 8678 6358 8730
rect 6358 8678 6404 8730
rect 6108 8676 6164 8678
rect 6188 8676 6244 8678
rect 6268 8676 6324 8678
rect 6348 8676 6404 8678
rect 3532 8186 3588 8188
rect 3612 8186 3668 8188
rect 3692 8186 3748 8188
rect 3772 8186 3828 8188
rect 3532 8134 3578 8186
rect 3578 8134 3588 8186
rect 3612 8134 3642 8186
rect 3642 8134 3654 8186
rect 3654 8134 3668 8186
rect 3692 8134 3706 8186
rect 3706 8134 3718 8186
rect 3718 8134 3748 8186
rect 3772 8134 3782 8186
rect 3782 8134 3828 8186
rect 3532 8132 3588 8134
rect 3612 8132 3668 8134
rect 3692 8132 3748 8134
rect 3772 8132 3828 8134
rect 6108 7642 6164 7644
rect 6188 7642 6244 7644
rect 6268 7642 6324 7644
rect 6348 7642 6404 7644
rect 6108 7590 6154 7642
rect 6154 7590 6164 7642
rect 6188 7590 6218 7642
rect 6218 7590 6230 7642
rect 6230 7590 6244 7642
rect 6268 7590 6282 7642
rect 6282 7590 6294 7642
rect 6294 7590 6324 7642
rect 6348 7590 6358 7642
rect 6358 7590 6404 7642
rect 6108 7588 6164 7590
rect 6188 7588 6244 7590
rect 6268 7588 6324 7590
rect 6348 7588 6404 7590
rect 3532 7098 3588 7100
rect 3612 7098 3668 7100
rect 3692 7098 3748 7100
rect 3772 7098 3828 7100
rect 3532 7046 3578 7098
rect 3578 7046 3588 7098
rect 3612 7046 3642 7098
rect 3642 7046 3654 7098
rect 3654 7046 3668 7098
rect 3692 7046 3706 7098
rect 3706 7046 3718 7098
rect 3718 7046 3748 7098
rect 3772 7046 3782 7098
rect 3782 7046 3828 7098
rect 3532 7044 3588 7046
rect 3612 7044 3668 7046
rect 3692 7044 3748 7046
rect 3772 7044 3828 7046
rect 6108 6554 6164 6556
rect 6188 6554 6244 6556
rect 6268 6554 6324 6556
rect 6348 6554 6404 6556
rect 6108 6502 6154 6554
rect 6154 6502 6164 6554
rect 6188 6502 6218 6554
rect 6218 6502 6230 6554
rect 6230 6502 6244 6554
rect 6268 6502 6282 6554
rect 6282 6502 6294 6554
rect 6294 6502 6324 6554
rect 6348 6502 6358 6554
rect 6358 6502 6404 6554
rect 6108 6500 6164 6502
rect 6188 6500 6244 6502
rect 6268 6500 6324 6502
rect 6348 6500 6404 6502
rect 3532 6010 3588 6012
rect 3612 6010 3668 6012
rect 3692 6010 3748 6012
rect 3772 6010 3828 6012
rect 3532 5958 3578 6010
rect 3578 5958 3588 6010
rect 3612 5958 3642 6010
rect 3642 5958 3654 6010
rect 3654 5958 3668 6010
rect 3692 5958 3706 6010
rect 3706 5958 3718 6010
rect 3718 5958 3748 6010
rect 3772 5958 3782 6010
rect 3782 5958 3828 6010
rect 3532 5956 3588 5958
rect 3612 5956 3668 5958
rect 3692 5956 3748 5958
rect 3772 5956 3828 5958
rect 6108 5466 6164 5468
rect 6188 5466 6244 5468
rect 6268 5466 6324 5468
rect 6348 5466 6404 5468
rect 6108 5414 6154 5466
rect 6154 5414 6164 5466
rect 6188 5414 6218 5466
rect 6218 5414 6230 5466
rect 6230 5414 6244 5466
rect 6268 5414 6282 5466
rect 6282 5414 6294 5466
rect 6294 5414 6324 5466
rect 6348 5414 6358 5466
rect 6358 5414 6404 5466
rect 6108 5412 6164 5414
rect 6188 5412 6244 5414
rect 6268 5412 6324 5414
rect 6348 5412 6404 5414
rect 8684 16890 8740 16892
rect 8764 16890 8820 16892
rect 8844 16890 8900 16892
rect 8924 16890 8980 16892
rect 8684 16838 8730 16890
rect 8730 16838 8740 16890
rect 8764 16838 8794 16890
rect 8794 16838 8806 16890
rect 8806 16838 8820 16890
rect 8844 16838 8858 16890
rect 8858 16838 8870 16890
rect 8870 16838 8900 16890
rect 8924 16838 8934 16890
rect 8934 16838 8980 16890
rect 8684 16836 8740 16838
rect 8764 16836 8820 16838
rect 8844 16836 8900 16838
rect 8924 16836 8980 16838
rect 13836 16890 13892 16892
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 13836 16838 13882 16890
rect 13882 16838 13892 16890
rect 13916 16838 13946 16890
rect 13946 16838 13958 16890
rect 13958 16838 13972 16890
rect 13996 16838 14010 16890
rect 14010 16838 14022 16890
rect 14022 16838 14052 16890
rect 14076 16838 14086 16890
rect 14086 16838 14132 16890
rect 13836 16836 13892 16838
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 11260 16346 11316 16348
rect 11340 16346 11396 16348
rect 11420 16346 11476 16348
rect 11500 16346 11556 16348
rect 11260 16294 11306 16346
rect 11306 16294 11316 16346
rect 11340 16294 11370 16346
rect 11370 16294 11382 16346
rect 11382 16294 11396 16346
rect 11420 16294 11434 16346
rect 11434 16294 11446 16346
rect 11446 16294 11476 16346
rect 11500 16294 11510 16346
rect 11510 16294 11556 16346
rect 11260 16292 11316 16294
rect 11340 16292 11396 16294
rect 11420 16292 11476 16294
rect 11500 16292 11556 16294
rect 8684 15802 8740 15804
rect 8764 15802 8820 15804
rect 8844 15802 8900 15804
rect 8924 15802 8980 15804
rect 8684 15750 8730 15802
rect 8730 15750 8740 15802
rect 8764 15750 8794 15802
rect 8794 15750 8806 15802
rect 8806 15750 8820 15802
rect 8844 15750 8858 15802
rect 8858 15750 8870 15802
rect 8870 15750 8900 15802
rect 8924 15750 8934 15802
rect 8934 15750 8980 15802
rect 8684 15748 8740 15750
rect 8764 15748 8820 15750
rect 8844 15748 8900 15750
rect 8924 15748 8980 15750
rect 13836 15802 13892 15804
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 13836 15750 13882 15802
rect 13882 15750 13892 15802
rect 13916 15750 13946 15802
rect 13946 15750 13958 15802
rect 13958 15750 13972 15802
rect 13996 15750 14010 15802
rect 14010 15750 14022 15802
rect 14022 15750 14052 15802
rect 14076 15750 14086 15802
rect 14086 15750 14132 15802
rect 13836 15748 13892 15750
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 8684 14714 8740 14716
rect 8764 14714 8820 14716
rect 8844 14714 8900 14716
rect 8924 14714 8980 14716
rect 8684 14662 8730 14714
rect 8730 14662 8740 14714
rect 8764 14662 8794 14714
rect 8794 14662 8806 14714
rect 8806 14662 8820 14714
rect 8844 14662 8858 14714
rect 8858 14662 8870 14714
rect 8870 14662 8900 14714
rect 8924 14662 8934 14714
rect 8934 14662 8980 14714
rect 8684 14660 8740 14662
rect 8764 14660 8820 14662
rect 8844 14660 8900 14662
rect 8924 14660 8980 14662
rect 8684 13626 8740 13628
rect 8764 13626 8820 13628
rect 8844 13626 8900 13628
rect 8924 13626 8980 13628
rect 8684 13574 8730 13626
rect 8730 13574 8740 13626
rect 8764 13574 8794 13626
rect 8794 13574 8806 13626
rect 8806 13574 8820 13626
rect 8844 13574 8858 13626
rect 8858 13574 8870 13626
rect 8870 13574 8900 13626
rect 8924 13574 8934 13626
rect 8934 13574 8980 13626
rect 8684 13572 8740 13574
rect 8764 13572 8820 13574
rect 8844 13572 8900 13574
rect 8924 13572 8980 13574
rect 8684 12538 8740 12540
rect 8764 12538 8820 12540
rect 8844 12538 8900 12540
rect 8924 12538 8980 12540
rect 8684 12486 8730 12538
rect 8730 12486 8740 12538
rect 8764 12486 8794 12538
rect 8794 12486 8806 12538
rect 8806 12486 8820 12538
rect 8844 12486 8858 12538
rect 8858 12486 8870 12538
rect 8870 12486 8900 12538
rect 8924 12486 8934 12538
rect 8934 12486 8980 12538
rect 8684 12484 8740 12486
rect 8764 12484 8820 12486
rect 8844 12484 8900 12486
rect 8924 12484 8980 12486
rect 8684 11450 8740 11452
rect 8764 11450 8820 11452
rect 8844 11450 8900 11452
rect 8924 11450 8980 11452
rect 8684 11398 8730 11450
rect 8730 11398 8740 11450
rect 8764 11398 8794 11450
rect 8794 11398 8806 11450
rect 8806 11398 8820 11450
rect 8844 11398 8858 11450
rect 8858 11398 8870 11450
rect 8870 11398 8900 11450
rect 8924 11398 8934 11450
rect 8934 11398 8980 11450
rect 8684 11396 8740 11398
rect 8764 11396 8820 11398
rect 8844 11396 8900 11398
rect 8924 11396 8980 11398
rect 8684 10362 8740 10364
rect 8764 10362 8820 10364
rect 8844 10362 8900 10364
rect 8924 10362 8980 10364
rect 8684 10310 8730 10362
rect 8730 10310 8740 10362
rect 8764 10310 8794 10362
rect 8794 10310 8806 10362
rect 8806 10310 8820 10362
rect 8844 10310 8858 10362
rect 8858 10310 8870 10362
rect 8870 10310 8900 10362
rect 8924 10310 8934 10362
rect 8934 10310 8980 10362
rect 8684 10308 8740 10310
rect 8764 10308 8820 10310
rect 8844 10308 8900 10310
rect 8924 10308 8980 10310
rect 8684 9274 8740 9276
rect 8764 9274 8820 9276
rect 8844 9274 8900 9276
rect 8924 9274 8980 9276
rect 8684 9222 8730 9274
rect 8730 9222 8740 9274
rect 8764 9222 8794 9274
rect 8794 9222 8806 9274
rect 8806 9222 8820 9274
rect 8844 9222 8858 9274
rect 8858 9222 8870 9274
rect 8870 9222 8900 9274
rect 8924 9222 8934 9274
rect 8934 9222 8980 9274
rect 8684 9220 8740 9222
rect 8764 9220 8820 9222
rect 8844 9220 8900 9222
rect 8924 9220 8980 9222
rect 8684 8186 8740 8188
rect 8764 8186 8820 8188
rect 8844 8186 8900 8188
rect 8924 8186 8980 8188
rect 8684 8134 8730 8186
rect 8730 8134 8740 8186
rect 8764 8134 8794 8186
rect 8794 8134 8806 8186
rect 8806 8134 8820 8186
rect 8844 8134 8858 8186
rect 8858 8134 8870 8186
rect 8870 8134 8900 8186
rect 8924 8134 8934 8186
rect 8934 8134 8980 8186
rect 8684 8132 8740 8134
rect 8764 8132 8820 8134
rect 8844 8132 8900 8134
rect 8924 8132 8980 8134
rect 8684 7098 8740 7100
rect 8764 7098 8820 7100
rect 8844 7098 8900 7100
rect 8924 7098 8980 7100
rect 8684 7046 8730 7098
rect 8730 7046 8740 7098
rect 8764 7046 8794 7098
rect 8794 7046 8806 7098
rect 8806 7046 8820 7098
rect 8844 7046 8858 7098
rect 8858 7046 8870 7098
rect 8870 7046 8900 7098
rect 8924 7046 8934 7098
rect 8934 7046 8980 7098
rect 8684 7044 8740 7046
rect 8764 7044 8820 7046
rect 8844 7044 8900 7046
rect 8924 7044 8980 7046
rect 8684 6010 8740 6012
rect 8764 6010 8820 6012
rect 8844 6010 8900 6012
rect 8924 6010 8980 6012
rect 8684 5958 8730 6010
rect 8730 5958 8740 6010
rect 8764 5958 8794 6010
rect 8794 5958 8806 6010
rect 8806 5958 8820 6010
rect 8844 5958 8858 6010
rect 8858 5958 8870 6010
rect 8870 5958 8900 6010
rect 8924 5958 8934 6010
rect 8934 5958 8980 6010
rect 8684 5956 8740 5958
rect 8764 5956 8820 5958
rect 8844 5956 8900 5958
rect 8924 5956 8980 5958
rect 3532 4922 3588 4924
rect 3612 4922 3668 4924
rect 3692 4922 3748 4924
rect 3772 4922 3828 4924
rect 3532 4870 3578 4922
rect 3578 4870 3588 4922
rect 3612 4870 3642 4922
rect 3642 4870 3654 4922
rect 3654 4870 3668 4922
rect 3692 4870 3706 4922
rect 3706 4870 3718 4922
rect 3718 4870 3748 4922
rect 3772 4870 3782 4922
rect 3782 4870 3828 4922
rect 3532 4868 3588 4870
rect 3612 4868 3668 4870
rect 3692 4868 3748 4870
rect 3772 4868 3828 4870
rect 6108 4378 6164 4380
rect 6188 4378 6244 4380
rect 6268 4378 6324 4380
rect 6348 4378 6404 4380
rect 6108 4326 6154 4378
rect 6154 4326 6164 4378
rect 6188 4326 6218 4378
rect 6218 4326 6230 4378
rect 6230 4326 6244 4378
rect 6268 4326 6282 4378
rect 6282 4326 6294 4378
rect 6294 4326 6324 4378
rect 6348 4326 6358 4378
rect 6358 4326 6404 4378
rect 6108 4324 6164 4326
rect 6188 4324 6244 4326
rect 6268 4324 6324 4326
rect 6348 4324 6404 4326
rect 3532 3834 3588 3836
rect 3612 3834 3668 3836
rect 3692 3834 3748 3836
rect 3772 3834 3828 3836
rect 3532 3782 3578 3834
rect 3578 3782 3588 3834
rect 3612 3782 3642 3834
rect 3642 3782 3654 3834
rect 3654 3782 3668 3834
rect 3692 3782 3706 3834
rect 3706 3782 3718 3834
rect 3718 3782 3748 3834
rect 3772 3782 3782 3834
rect 3782 3782 3828 3834
rect 3532 3780 3588 3782
rect 3612 3780 3668 3782
rect 3692 3780 3748 3782
rect 3772 3780 3828 3782
rect 6108 3290 6164 3292
rect 6188 3290 6244 3292
rect 6268 3290 6324 3292
rect 6348 3290 6404 3292
rect 6108 3238 6154 3290
rect 6154 3238 6164 3290
rect 6188 3238 6218 3290
rect 6218 3238 6230 3290
rect 6230 3238 6244 3290
rect 6268 3238 6282 3290
rect 6282 3238 6294 3290
rect 6294 3238 6324 3290
rect 6348 3238 6358 3290
rect 6358 3238 6404 3290
rect 6108 3236 6164 3238
rect 6188 3236 6244 3238
rect 6268 3236 6324 3238
rect 6348 3236 6404 3238
rect 3532 2746 3588 2748
rect 3612 2746 3668 2748
rect 3692 2746 3748 2748
rect 3772 2746 3828 2748
rect 3532 2694 3578 2746
rect 3578 2694 3588 2746
rect 3612 2694 3642 2746
rect 3642 2694 3654 2746
rect 3654 2694 3668 2746
rect 3692 2694 3706 2746
rect 3706 2694 3718 2746
rect 3718 2694 3748 2746
rect 3772 2694 3782 2746
rect 3782 2694 3828 2746
rect 3532 2692 3588 2694
rect 3612 2692 3668 2694
rect 3692 2692 3748 2694
rect 3772 2692 3828 2694
rect 8684 4922 8740 4924
rect 8764 4922 8820 4924
rect 8844 4922 8900 4924
rect 8924 4922 8980 4924
rect 8684 4870 8730 4922
rect 8730 4870 8740 4922
rect 8764 4870 8794 4922
rect 8794 4870 8806 4922
rect 8806 4870 8820 4922
rect 8844 4870 8858 4922
rect 8858 4870 8870 4922
rect 8870 4870 8900 4922
rect 8924 4870 8934 4922
rect 8934 4870 8980 4922
rect 8684 4868 8740 4870
rect 8764 4868 8820 4870
rect 8844 4868 8900 4870
rect 8924 4868 8980 4870
rect 11260 15258 11316 15260
rect 11340 15258 11396 15260
rect 11420 15258 11476 15260
rect 11500 15258 11556 15260
rect 11260 15206 11306 15258
rect 11306 15206 11316 15258
rect 11340 15206 11370 15258
rect 11370 15206 11382 15258
rect 11382 15206 11396 15258
rect 11420 15206 11434 15258
rect 11434 15206 11446 15258
rect 11446 15206 11476 15258
rect 11500 15206 11510 15258
rect 11510 15206 11556 15258
rect 11260 15204 11316 15206
rect 11340 15204 11396 15206
rect 11420 15204 11476 15206
rect 11500 15204 11556 15206
rect 13836 14714 13892 14716
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 13836 14662 13882 14714
rect 13882 14662 13892 14714
rect 13916 14662 13946 14714
rect 13946 14662 13958 14714
rect 13958 14662 13972 14714
rect 13996 14662 14010 14714
rect 14010 14662 14022 14714
rect 14022 14662 14052 14714
rect 14076 14662 14086 14714
rect 14086 14662 14132 14714
rect 13836 14660 13892 14662
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 11260 14170 11316 14172
rect 11340 14170 11396 14172
rect 11420 14170 11476 14172
rect 11500 14170 11556 14172
rect 11260 14118 11306 14170
rect 11306 14118 11316 14170
rect 11340 14118 11370 14170
rect 11370 14118 11382 14170
rect 11382 14118 11396 14170
rect 11420 14118 11434 14170
rect 11434 14118 11446 14170
rect 11446 14118 11476 14170
rect 11500 14118 11510 14170
rect 11510 14118 11556 14170
rect 11260 14116 11316 14118
rect 11340 14116 11396 14118
rect 11420 14116 11476 14118
rect 11500 14116 11556 14118
rect 13836 13626 13892 13628
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 13836 13574 13882 13626
rect 13882 13574 13892 13626
rect 13916 13574 13946 13626
rect 13946 13574 13958 13626
rect 13958 13574 13972 13626
rect 13996 13574 14010 13626
rect 14010 13574 14022 13626
rect 14022 13574 14052 13626
rect 14076 13574 14086 13626
rect 14086 13574 14132 13626
rect 13836 13572 13892 13574
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 11260 13082 11316 13084
rect 11340 13082 11396 13084
rect 11420 13082 11476 13084
rect 11500 13082 11556 13084
rect 11260 13030 11306 13082
rect 11306 13030 11316 13082
rect 11340 13030 11370 13082
rect 11370 13030 11382 13082
rect 11382 13030 11396 13082
rect 11420 13030 11434 13082
rect 11434 13030 11446 13082
rect 11446 13030 11476 13082
rect 11500 13030 11510 13082
rect 11510 13030 11556 13082
rect 11260 13028 11316 13030
rect 11340 13028 11396 13030
rect 11420 13028 11476 13030
rect 11500 13028 11556 13030
rect 13836 12538 13892 12540
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 13836 12486 13882 12538
rect 13882 12486 13892 12538
rect 13916 12486 13946 12538
rect 13946 12486 13958 12538
rect 13958 12486 13972 12538
rect 13996 12486 14010 12538
rect 14010 12486 14022 12538
rect 14022 12486 14052 12538
rect 14076 12486 14086 12538
rect 14086 12486 14132 12538
rect 13836 12484 13892 12486
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 11260 11994 11316 11996
rect 11340 11994 11396 11996
rect 11420 11994 11476 11996
rect 11500 11994 11556 11996
rect 11260 11942 11306 11994
rect 11306 11942 11316 11994
rect 11340 11942 11370 11994
rect 11370 11942 11382 11994
rect 11382 11942 11396 11994
rect 11420 11942 11434 11994
rect 11434 11942 11446 11994
rect 11446 11942 11476 11994
rect 11500 11942 11510 11994
rect 11510 11942 11556 11994
rect 11260 11940 11316 11942
rect 11340 11940 11396 11942
rect 11420 11940 11476 11942
rect 11500 11940 11556 11942
rect 13836 11450 13892 11452
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 13836 11398 13882 11450
rect 13882 11398 13892 11450
rect 13916 11398 13946 11450
rect 13946 11398 13958 11450
rect 13958 11398 13972 11450
rect 13996 11398 14010 11450
rect 14010 11398 14022 11450
rect 14022 11398 14052 11450
rect 14076 11398 14086 11450
rect 14086 11398 14132 11450
rect 13836 11396 13892 11398
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 11260 10906 11316 10908
rect 11340 10906 11396 10908
rect 11420 10906 11476 10908
rect 11500 10906 11556 10908
rect 11260 10854 11306 10906
rect 11306 10854 11316 10906
rect 11340 10854 11370 10906
rect 11370 10854 11382 10906
rect 11382 10854 11396 10906
rect 11420 10854 11434 10906
rect 11434 10854 11446 10906
rect 11446 10854 11476 10906
rect 11500 10854 11510 10906
rect 11510 10854 11556 10906
rect 11260 10852 11316 10854
rect 11340 10852 11396 10854
rect 11420 10852 11476 10854
rect 11500 10852 11556 10854
rect 13836 10362 13892 10364
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 13836 10310 13882 10362
rect 13882 10310 13892 10362
rect 13916 10310 13946 10362
rect 13946 10310 13958 10362
rect 13958 10310 13972 10362
rect 13996 10310 14010 10362
rect 14010 10310 14022 10362
rect 14022 10310 14052 10362
rect 14076 10310 14086 10362
rect 14086 10310 14132 10362
rect 13836 10308 13892 10310
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 11260 9818 11316 9820
rect 11340 9818 11396 9820
rect 11420 9818 11476 9820
rect 11500 9818 11556 9820
rect 11260 9766 11306 9818
rect 11306 9766 11316 9818
rect 11340 9766 11370 9818
rect 11370 9766 11382 9818
rect 11382 9766 11396 9818
rect 11420 9766 11434 9818
rect 11434 9766 11446 9818
rect 11446 9766 11476 9818
rect 11500 9766 11510 9818
rect 11510 9766 11556 9818
rect 11260 9764 11316 9766
rect 11340 9764 11396 9766
rect 11420 9764 11476 9766
rect 11500 9764 11556 9766
rect 13836 9274 13892 9276
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 13836 9222 13882 9274
rect 13882 9222 13892 9274
rect 13916 9222 13946 9274
rect 13946 9222 13958 9274
rect 13958 9222 13972 9274
rect 13996 9222 14010 9274
rect 14010 9222 14022 9274
rect 14022 9222 14052 9274
rect 14076 9222 14086 9274
rect 14086 9222 14132 9274
rect 13836 9220 13892 9222
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 11260 8730 11316 8732
rect 11340 8730 11396 8732
rect 11420 8730 11476 8732
rect 11500 8730 11556 8732
rect 11260 8678 11306 8730
rect 11306 8678 11316 8730
rect 11340 8678 11370 8730
rect 11370 8678 11382 8730
rect 11382 8678 11396 8730
rect 11420 8678 11434 8730
rect 11434 8678 11446 8730
rect 11446 8678 11476 8730
rect 11500 8678 11510 8730
rect 11510 8678 11556 8730
rect 11260 8676 11316 8678
rect 11340 8676 11396 8678
rect 11420 8676 11476 8678
rect 11500 8676 11556 8678
rect 13836 8186 13892 8188
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 13836 8134 13882 8186
rect 13882 8134 13892 8186
rect 13916 8134 13946 8186
rect 13946 8134 13958 8186
rect 13958 8134 13972 8186
rect 13996 8134 14010 8186
rect 14010 8134 14022 8186
rect 14022 8134 14052 8186
rect 14076 8134 14086 8186
rect 14086 8134 14132 8186
rect 13836 8132 13892 8134
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 11260 7642 11316 7644
rect 11340 7642 11396 7644
rect 11420 7642 11476 7644
rect 11500 7642 11556 7644
rect 11260 7590 11306 7642
rect 11306 7590 11316 7642
rect 11340 7590 11370 7642
rect 11370 7590 11382 7642
rect 11382 7590 11396 7642
rect 11420 7590 11434 7642
rect 11434 7590 11446 7642
rect 11446 7590 11476 7642
rect 11500 7590 11510 7642
rect 11510 7590 11556 7642
rect 11260 7588 11316 7590
rect 11340 7588 11396 7590
rect 11420 7588 11476 7590
rect 11500 7588 11556 7590
rect 13836 7098 13892 7100
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 13836 7046 13882 7098
rect 13882 7046 13892 7098
rect 13916 7046 13946 7098
rect 13946 7046 13958 7098
rect 13958 7046 13972 7098
rect 13996 7046 14010 7098
rect 14010 7046 14022 7098
rect 14022 7046 14052 7098
rect 14076 7046 14086 7098
rect 14086 7046 14132 7098
rect 13836 7044 13892 7046
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 11260 6554 11316 6556
rect 11340 6554 11396 6556
rect 11420 6554 11476 6556
rect 11500 6554 11556 6556
rect 11260 6502 11306 6554
rect 11306 6502 11316 6554
rect 11340 6502 11370 6554
rect 11370 6502 11382 6554
rect 11382 6502 11396 6554
rect 11420 6502 11434 6554
rect 11434 6502 11446 6554
rect 11446 6502 11476 6554
rect 11500 6502 11510 6554
rect 11510 6502 11556 6554
rect 11260 6500 11316 6502
rect 11340 6500 11396 6502
rect 11420 6500 11476 6502
rect 11500 6500 11556 6502
rect 13836 6010 13892 6012
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 13836 5958 13882 6010
rect 13882 5958 13892 6010
rect 13916 5958 13946 6010
rect 13946 5958 13958 6010
rect 13958 5958 13972 6010
rect 13996 5958 14010 6010
rect 14010 5958 14022 6010
rect 14022 5958 14052 6010
rect 14076 5958 14086 6010
rect 14086 5958 14132 6010
rect 13836 5956 13892 5958
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 11260 5466 11316 5468
rect 11340 5466 11396 5468
rect 11420 5466 11476 5468
rect 11500 5466 11556 5468
rect 11260 5414 11306 5466
rect 11306 5414 11316 5466
rect 11340 5414 11370 5466
rect 11370 5414 11382 5466
rect 11382 5414 11396 5466
rect 11420 5414 11434 5466
rect 11434 5414 11446 5466
rect 11446 5414 11476 5466
rect 11500 5414 11510 5466
rect 11510 5414 11556 5466
rect 11260 5412 11316 5414
rect 11340 5412 11396 5414
rect 11420 5412 11476 5414
rect 11500 5412 11556 5414
rect 8684 3834 8740 3836
rect 8764 3834 8820 3836
rect 8844 3834 8900 3836
rect 8924 3834 8980 3836
rect 8684 3782 8730 3834
rect 8730 3782 8740 3834
rect 8764 3782 8794 3834
rect 8794 3782 8806 3834
rect 8806 3782 8820 3834
rect 8844 3782 8858 3834
rect 8858 3782 8870 3834
rect 8870 3782 8900 3834
rect 8924 3782 8934 3834
rect 8934 3782 8980 3834
rect 8684 3780 8740 3782
rect 8764 3780 8820 3782
rect 8844 3780 8900 3782
rect 8924 3780 8980 3782
rect 8684 2746 8740 2748
rect 8764 2746 8820 2748
rect 8844 2746 8900 2748
rect 8924 2746 8980 2748
rect 8684 2694 8730 2746
rect 8730 2694 8740 2746
rect 8764 2694 8794 2746
rect 8794 2694 8806 2746
rect 8806 2694 8820 2746
rect 8844 2694 8858 2746
rect 8858 2694 8870 2746
rect 8870 2694 8900 2746
rect 8924 2694 8934 2746
rect 8934 2694 8980 2746
rect 8684 2692 8740 2694
rect 8764 2692 8820 2694
rect 8844 2692 8900 2694
rect 8924 2692 8980 2694
rect 13836 4922 13892 4924
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 13836 4870 13882 4922
rect 13882 4870 13892 4922
rect 13916 4870 13946 4922
rect 13946 4870 13958 4922
rect 13958 4870 13972 4922
rect 13996 4870 14010 4922
rect 14010 4870 14022 4922
rect 14022 4870 14052 4922
rect 14076 4870 14086 4922
rect 14086 4870 14132 4922
rect 13836 4868 13892 4870
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 11260 4378 11316 4380
rect 11340 4378 11396 4380
rect 11420 4378 11476 4380
rect 11500 4378 11556 4380
rect 11260 4326 11306 4378
rect 11306 4326 11316 4378
rect 11340 4326 11370 4378
rect 11370 4326 11382 4378
rect 11382 4326 11396 4378
rect 11420 4326 11434 4378
rect 11434 4326 11446 4378
rect 11446 4326 11476 4378
rect 11500 4326 11510 4378
rect 11510 4326 11556 4378
rect 11260 4324 11316 4326
rect 11340 4324 11396 4326
rect 11420 4324 11476 4326
rect 11500 4324 11556 4326
rect 11260 3290 11316 3292
rect 11340 3290 11396 3292
rect 11420 3290 11476 3292
rect 11500 3290 11556 3292
rect 11260 3238 11306 3290
rect 11306 3238 11316 3290
rect 11340 3238 11370 3290
rect 11370 3238 11382 3290
rect 11382 3238 11396 3290
rect 11420 3238 11434 3290
rect 11434 3238 11446 3290
rect 11446 3238 11476 3290
rect 11500 3238 11510 3290
rect 11510 3238 11556 3290
rect 11260 3236 11316 3238
rect 11340 3236 11396 3238
rect 11420 3236 11476 3238
rect 11500 3236 11556 3238
rect 13836 3834 13892 3836
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 13836 3782 13882 3834
rect 13882 3782 13892 3834
rect 13916 3782 13946 3834
rect 13946 3782 13958 3834
rect 13958 3782 13972 3834
rect 13996 3782 14010 3834
rect 14010 3782 14022 3834
rect 14022 3782 14052 3834
rect 14076 3782 14086 3834
rect 14086 3782 14132 3834
rect 13836 3780 13892 3782
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 13836 2746 13892 2748
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 13836 2694 13882 2746
rect 13882 2694 13892 2746
rect 13916 2694 13946 2746
rect 13946 2694 13958 2746
rect 13958 2694 13972 2746
rect 13996 2694 14010 2746
rect 14010 2694 14022 2746
rect 14022 2694 14052 2746
rect 14076 2694 14086 2746
rect 14086 2694 14132 2746
rect 13836 2692 13892 2694
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 6108 2202 6164 2204
rect 6188 2202 6244 2204
rect 6268 2202 6324 2204
rect 6348 2202 6404 2204
rect 6108 2150 6154 2202
rect 6154 2150 6164 2202
rect 6188 2150 6218 2202
rect 6218 2150 6230 2202
rect 6230 2150 6244 2202
rect 6268 2150 6282 2202
rect 6282 2150 6294 2202
rect 6294 2150 6324 2202
rect 6348 2150 6358 2202
rect 6358 2150 6404 2202
rect 6108 2148 6164 2150
rect 6188 2148 6244 2150
rect 6268 2148 6324 2150
rect 6348 2148 6404 2150
rect 11260 2202 11316 2204
rect 11340 2202 11396 2204
rect 11420 2202 11476 2204
rect 11500 2202 11556 2204
rect 11260 2150 11306 2202
rect 11306 2150 11316 2202
rect 11340 2150 11370 2202
rect 11370 2150 11382 2202
rect 11382 2150 11396 2202
rect 11420 2150 11434 2202
rect 11434 2150 11446 2202
rect 11446 2150 11476 2202
rect 11500 2150 11510 2202
rect 11510 2150 11556 2202
rect 11260 2148 11316 2150
rect 11340 2148 11396 2150
rect 11420 2148 11476 2150
rect 11500 2148 11556 2150
<< metal3 >>
rect 6096 17440 6416 17441
rect 6096 17376 6104 17440
rect 6168 17376 6184 17440
rect 6248 17376 6264 17440
rect 6328 17376 6344 17440
rect 6408 17376 6416 17440
rect 6096 17375 6416 17376
rect 11248 17440 11568 17441
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 17375 11568 17376
rect 3520 16896 3840 16897
rect 3520 16832 3528 16896
rect 3592 16832 3608 16896
rect 3672 16832 3688 16896
rect 3752 16832 3768 16896
rect 3832 16832 3840 16896
rect 3520 16831 3840 16832
rect 8672 16896 8992 16897
rect 8672 16832 8680 16896
rect 8744 16832 8760 16896
rect 8824 16832 8840 16896
rect 8904 16832 8920 16896
rect 8984 16832 8992 16896
rect 8672 16831 8992 16832
rect 13824 16896 14144 16897
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 13824 16831 14144 16832
rect 6096 16352 6416 16353
rect 6096 16288 6104 16352
rect 6168 16288 6184 16352
rect 6248 16288 6264 16352
rect 6328 16288 6344 16352
rect 6408 16288 6416 16352
rect 6096 16287 6416 16288
rect 11248 16352 11568 16353
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 16287 11568 16288
rect 3520 15808 3840 15809
rect 3520 15744 3528 15808
rect 3592 15744 3608 15808
rect 3672 15744 3688 15808
rect 3752 15744 3768 15808
rect 3832 15744 3840 15808
rect 3520 15743 3840 15744
rect 8672 15808 8992 15809
rect 8672 15744 8680 15808
rect 8744 15744 8760 15808
rect 8824 15744 8840 15808
rect 8904 15744 8920 15808
rect 8984 15744 8992 15808
rect 8672 15743 8992 15744
rect 13824 15808 14144 15809
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 15743 14144 15744
rect 6096 15264 6416 15265
rect 6096 15200 6104 15264
rect 6168 15200 6184 15264
rect 6248 15200 6264 15264
rect 6328 15200 6344 15264
rect 6408 15200 6416 15264
rect 6096 15199 6416 15200
rect 11248 15264 11568 15265
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 15199 11568 15200
rect 3520 14720 3840 14721
rect 3520 14656 3528 14720
rect 3592 14656 3608 14720
rect 3672 14656 3688 14720
rect 3752 14656 3768 14720
rect 3832 14656 3840 14720
rect 3520 14655 3840 14656
rect 8672 14720 8992 14721
rect 8672 14656 8680 14720
rect 8744 14656 8760 14720
rect 8824 14656 8840 14720
rect 8904 14656 8920 14720
rect 8984 14656 8992 14720
rect 8672 14655 8992 14656
rect 13824 14720 14144 14721
rect 13824 14656 13832 14720
rect 13896 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14144 14720
rect 13824 14655 14144 14656
rect 6096 14176 6416 14177
rect 6096 14112 6104 14176
rect 6168 14112 6184 14176
rect 6248 14112 6264 14176
rect 6328 14112 6344 14176
rect 6408 14112 6416 14176
rect 6096 14111 6416 14112
rect 11248 14176 11568 14177
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 14111 11568 14112
rect 3520 13632 3840 13633
rect 3520 13568 3528 13632
rect 3592 13568 3608 13632
rect 3672 13568 3688 13632
rect 3752 13568 3768 13632
rect 3832 13568 3840 13632
rect 3520 13567 3840 13568
rect 8672 13632 8992 13633
rect 8672 13568 8680 13632
rect 8744 13568 8760 13632
rect 8824 13568 8840 13632
rect 8904 13568 8920 13632
rect 8984 13568 8992 13632
rect 8672 13567 8992 13568
rect 13824 13632 14144 13633
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 13567 14144 13568
rect 6096 13088 6416 13089
rect 6096 13024 6104 13088
rect 6168 13024 6184 13088
rect 6248 13024 6264 13088
rect 6328 13024 6344 13088
rect 6408 13024 6416 13088
rect 6096 13023 6416 13024
rect 11248 13088 11568 13089
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 13023 11568 13024
rect 3520 12544 3840 12545
rect 3520 12480 3528 12544
rect 3592 12480 3608 12544
rect 3672 12480 3688 12544
rect 3752 12480 3768 12544
rect 3832 12480 3840 12544
rect 3520 12479 3840 12480
rect 8672 12544 8992 12545
rect 8672 12480 8680 12544
rect 8744 12480 8760 12544
rect 8824 12480 8840 12544
rect 8904 12480 8920 12544
rect 8984 12480 8992 12544
rect 8672 12479 8992 12480
rect 13824 12544 14144 12545
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 12479 14144 12480
rect 6096 12000 6416 12001
rect 6096 11936 6104 12000
rect 6168 11936 6184 12000
rect 6248 11936 6264 12000
rect 6328 11936 6344 12000
rect 6408 11936 6416 12000
rect 6096 11935 6416 11936
rect 11248 12000 11568 12001
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 11935 11568 11936
rect 3520 11456 3840 11457
rect 3520 11392 3528 11456
rect 3592 11392 3608 11456
rect 3672 11392 3688 11456
rect 3752 11392 3768 11456
rect 3832 11392 3840 11456
rect 3520 11391 3840 11392
rect 8672 11456 8992 11457
rect 8672 11392 8680 11456
rect 8744 11392 8760 11456
rect 8824 11392 8840 11456
rect 8904 11392 8920 11456
rect 8984 11392 8992 11456
rect 8672 11391 8992 11392
rect 13824 11456 14144 11457
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 11391 14144 11392
rect 6096 10912 6416 10913
rect 6096 10848 6104 10912
rect 6168 10848 6184 10912
rect 6248 10848 6264 10912
rect 6328 10848 6344 10912
rect 6408 10848 6416 10912
rect 6096 10847 6416 10848
rect 11248 10912 11568 10913
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 10847 11568 10848
rect 3520 10368 3840 10369
rect 3520 10304 3528 10368
rect 3592 10304 3608 10368
rect 3672 10304 3688 10368
rect 3752 10304 3768 10368
rect 3832 10304 3840 10368
rect 3520 10303 3840 10304
rect 8672 10368 8992 10369
rect 8672 10304 8680 10368
rect 8744 10304 8760 10368
rect 8824 10304 8840 10368
rect 8904 10304 8920 10368
rect 8984 10304 8992 10368
rect 8672 10303 8992 10304
rect 13824 10368 14144 10369
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 10303 14144 10304
rect 6096 9824 6416 9825
rect 6096 9760 6104 9824
rect 6168 9760 6184 9824
rect 6248 9760 6264 9824
rect 6328 9760 6344 9824
rect 6408 9760 6416 9824
rect 6096 9759 6416 9760
rect 11248 9824 11568 9825
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 9759 11568 9760
rect 3520 9280 3840 9281
rect 3520 9216 3528 9280
rect 3592 9216 3608 9280
rect 3672 9216 3688 9280
rect 3752 9216 3768 9280
rect 3832 9216 3840 9280
rect 3520 9215 3840 9216
rect 8672 9280 8992 9281
rect 8672 9216 8680 9280
rect 8744 9216 8760 9280
rect 8824 9216 8840 9280
rect 8904 9216 8920 9280
rect 8984 9216 8992 9280
rect 8672 9215 8992 9216
rect 13824 9280 14144 9281
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 9215 14144 9216
rect 6096 8736 6416 8737
rect 6096 8672 6104 8736
rect 6168 8672 6184 8736
rect 6248 8672 6264 8736
rect 6328 8672 6344 8736
rect 6408 8672 6416 8736
rect 6096 8671 6416 8672
rect 11248 8736 11568 8737
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 8671 11568 8672
rect 3520 8192 3840 8193
rect 3520 8128 3528 8192
rect 3592 8128 3608 8192
rect 3672 8128 3688 8192
rect 3752 8128 3768 8192
rect 3832 8128 3840 8192
rect 3520 8127 3840 8128
rect 8672 8192 8992 8193
rect 8672 8128 8680 8192
rect 8744 8128 8760 8192
rect 8824 8128 8840 8192
rect 8904 8128 8920 8192
rect 8984 8128 8992 8192
rect 8672 8127 8992 8128
rect 13824 8192 14144 8193
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 8127 14144 8128
rect 6096 7648 6416 7649
rect 6096 7584 6104 7648
rect 6168 7584 6184 7648
rect 6248 7584 6264 7648
rect 6328 7584 6344 7648
rect 6408 7584 6416 7648
rect 6096 7583 6416 7584
rect 11248 7648 11568 7649
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 7583 11568 7584
rect 3520 7104 3840 7105
rect 3520 7040 3528 7104
rect 3592 7040 3608 7104
rect 3672 7040 3688 7104
rect 3752 7040 3768 7104
rect 3832 7040 3840 7104
rect 3520 7039 3840 7040
rect 8672 7104 8992 7105
rect 8672 7040 8680 7104
rect 8744 7040 8760 7104
rect 8824 7040 8840 7104
rect 8904 7040 8920 7104
rect 8984 7040 8992 7104
rect 8672 7039 8992 7040
rect 13824 7104 14144 7105
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 7039 14144 7040
rect 6096 6560 6416 6561
rect 6096 6496 6104 6560
rect 6168 6496 6184 6560
rect 6248 6496 6264 6560
rect 6328 6496 6344 6560
rect 6408 6496 6416 6560
rect 6096 6495 6416 6496
rect 11248 6560 11568 6561
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 6495 11568 6496
rect 3520 6016 3840 6017
rect 3520 5952 3528 6016
rect 3592 5952 3608 6016
rect 3672 5952 3688 6016
rect 3752 5952 3768 6016
rect 3832 5952 3840 6016
rect 3520 5951 3840 5952
rect 8672 6016 8992 6017
rect 8672 5952 8680 6016
rect 8744 5952 8760 6016
rect 8824 5952 8840 6016
rect 8904 5952 8920 6016
rect 8984 5952 8992 6016
rect 8672 5951 8992 5952
rect 13824 6016 14144 6017
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 13824 5951 14144 5952
rect 6096 5472 6416 5473
rect 6096 5408 6104 5472
rect 6168 5408 6184 5472
rect 6248 5408 6264 5472
rect 6328 5408 6344 5472
rect 6408 5408 6416 5472
rect 6096 5407 6416 5408
rect 11248 5472 11568 5473
rect 11248 5408 11256 5472
rect 11320 5408 11336 5472
rect 11400 5408 11416 5472
rect 11480 5408 11496 5472
rect 11560 5408 11568 5472
rect 11248 5407 11568 5408
rect 3520 4928 3840 4929
rect 3520 4864 3528 4928
rect 3592 4864 3608 4928
rect 3672 4864 3688 4928
rect 3752 4864 3768 4928
rect 3832 4864 3840 4928
rect 3520 4863 3840 4864
rect 8672 4928 8992 4929
rect 8672 4864 8680 4928
rect 8744 4864 8760 4928
rect 8824 4864 8840 4928
rect 8904 4864 8920 4928
rect 8984 4864 8992 4928
rect 8672 4863 8992 4864
rect 13824 4928 14144 4929
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 4863 14144 4864
rect 6096 4384 6416 4385
rect 6096 4320 6104 4384
rect 6168 4320 6184 4384
rect 6248 4320 6264 4384
rect 6328 4320 6344 4384
rect 6408 4320 6416 4384
rect 6096 4319 6416 4320
rect 11248 4384 11568 4385
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 4319 11568 4320
rect 3520 3840 3840 3841
rect 3520 3776 3528 3840
rect 3592 3776 3608 3840
rect 3672 3776 3688 3840
rect 3752 3776 3768 3840
rect 3832 3776 3840 3840
rect 3520 3775 3840 3776
rect 8672 3840 8992 3841
rect 8672 3776 8680 3840
rect 8744 3776 8760 3840
rect 8824 3776 8840 3840
rect 8904 3776 8920 3840
rect 8984 3776 8992 3840
rect 8672 3775 8992 3776
rect 13824 3840 14144 3841
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 3775 14144 3776
rect 6096 3296 6416 3297
rect 6096 3232 6104 3296
rect 6168 3232 6184 3296
rect 6248 3232 6264 3296
rect 6328 3232 6344 3296
rect 6408 3232 6416 3296
rect 6096 3231 6416 3232
rect 11248 3296 11568 3297
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 3231 11568 3232
rect 3520 2752 3840 2753
rect 3520 2688 3528 2752
rect 3592 2688 3608 2752
rect 3672 2688 3688 2752
rect 3752 2688 3768 2752
rect 3832 2688 3840 2752
rect 3520 2687 3840 2688
rect 8672 2752 8992 2753
rect 8672 2688 8680 2752
rect 8744 2688 8760 2752
rect 8824 2688 8840 2752
rect 8904 2688 8920 2752
rect 8984 2688 8992 2752
rect 8672 2687 8992 2688
rect 13824 2752 14144 2753
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 2687 14144 2688
rect 6096 2208 6416 2209
rect 6096 2144 6104 2208
rect 6168 2144 6184 2208
rect 6248 2144 6264 2208
rect 6328 2144 6344 2208
rect 6408 2144 6416 2208
rect 6096 2143 6416 2144
rect 11248 2208 11568 2209
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2143 11568 2144
<< via3 >>
rect 6104 17436 6168 17440
rect 6104 17380 6108 17436
rect 6108 17380 6164 17436
rect 6164 17380 6168 17436
rect 6104 17376 6168 17380
rect 6184 17436 6248 17440
rect 6184 17380 6188 17436
rect 6188 17380 6244 17436
rect 6244 17380 6248 17436
rect 6184 17376 6248 17380
rect 6264 17436 6328 17440
rect 6264 17380 6268 17436
rect 6268 17380 6324 17436
rect 6324 17380 6328 17436
rect 6264 17376 6328 17380
rect 6344 17436 6408 17440
rect 6344 17380 6348 17436
rect 6348 17380 6404 17436
rect 6404 17380 6408 17436
rect 6344 17376 6408 17380
rect 11256 17436 11320 17440
rect 11256 17380 11260 17436
rect 11260 17380 11316 17436
rect 11316 17380 11320 17436
rect 11256 17376 11320 17380
rect 11336 17436 11400 17440
rect 11336 17380 11340 17436
rect 11340 17380 11396 17436
rect 11396 17380 11400 17436
rect 11336 17376 11400 17380
rect 11416 17436 11480 17440
rect 11416 17380 11420 17436
rect 11420 17380 11476 17436
rect 11476 17380 11480 17436
rect 11416 17376 11480 17380
rect 11496 17436 11560 17440
rect 11496 17380 11500 17436
rect 11500 17380 11556 17436
rect 11556 17380 11560 17436
rect 11496 17376 11560 17380
rect 3528 16892 3592 16896
rect 3528 16836 3532 16892
rect 3532 16836 3588 16892
rect 3588 16836 3592 16892
rect 3528 16832 3592 16836
rect 3608 16892 3672 16896
rect 3608 16836 3612 16892
rect 3612 16836 3668 16892
rect 3668 16836 3672 16892
rect 3608 16832 3672 16836
rect 3688 16892 3752 16896
rect 3688 16836 3692 16892
rect 3692 16836 3748 16892
rect 3748 16836 3752 16892
rect 3688 16832 3752 16836
rect 3768 16892 3832 16896
rect 3768 16836 3772 16892
rect 3772 16836 3828 16892
rect 3828 16836 3832 16892
rect 3768 16832 3832 16836
rect 8680 16892 8744 16896
rect 8680 16836 8684 16892
rect 8684 16836 8740 16892
rect 8740 16836 8744 16892
rect 8680 16832 8744 16836
rect 8760 16892 8824 16896
rect 8760 16836 8764 16892
rect 8764 16836 8820 16892
rect 8820 16836 8824 16892
rect 8760 16832 8824 16836
rect 8840 16892 8904 16896
rect 8840 16836 8844 16892
rect 8844 16836 8900 16892
rect 8900 16836 8904 16892
rect 8840 16832 8904 16836
rect 8920 16892 8984 16896
rect 8920 16836 8924 16892
rect 8924 16836 8980 16892
rect 8980 16836 8984 16892
rect 8920 16832 8984 16836
rect 13832 16892 13896 16896
rect 13832 16836 13836 16892
rect 13836 16836 13892 16892
rect 13892 16836 13896 16892
rect 13832 16832 13896 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 6104 16348 6168 16352
rect 6104 16292 6108 16348
rect 6108 16292 6164 16348
rect 6164 16292 6168 16348
rect 6104 16288 6168 16292
rect 6184 16348 6248 16352
rect 6184 16292 6188 16348
rect 6188 16292 6244 16348
rect 6244 16292 6248 16348
rect 6184 16288 6248 16292
rect 6264 16348 6328 16352
rect 6264 16292 6268 16348
rect 6268 16292 6324 16348
rect 6324 16292 6328 16348
rect 6264 16288 6328 16292
rect 6344 16348 6408 16352
rect 6344 16292 6348 16348
rect 6348 16292 6404 16348
rect 6404 16292 6408 16348
rect 6344 16288 6408 16292
rect 11256 16348 11320 16352
rect 11256 16292 11260 16348
rect 11260 16292 11316 16348
rect 11316 16292 11320 16348
rect 11256 16288 11320 16292
rect 11336 16348 11400 16352
rect 11336 16292 11340 16348
rect 11340 16292 11396 16348
rect 11396 16292 11400 16348
rect 11336 16288 11400 16292
rect 11416 16348 11480 16352
rect 11416 16292 11420 16348
rect 11420 16292 11476 16348
rect 11476 16292 11480 16348
rect 11416 16288 11480 16292
rect 11496 16348 11560 16352
rect 11496 16292 11500 16348
rect 11500 16292 11556 16348
rect 11556 16292 11560 16348
rect 11496 16288 11560 16292
rect 3528 15804 3592 15808
rect 3528 15748 3532 15804
rect 3532 15748 3588 15804
rect 3588 15748 3592 15804
rect 3528 15744 3592 15748
rect 3608 15804 3672 15808
rect 3608 15748 3612 15804
rect 3612 15748 3668 15804
rect 3668 15748 3672 15804
rect 3608 15744 3672 15748
rect 3688 15804 3752 15808
rect 3688 15748 3692 15804
rect 3692 15748 3748 15804
rect 3748 15748 3752 15804
rect 3688 15744 3752 15748
rect 3768 15804 3832 15808
rect 3768 15748 3772 15804
rect 3772 15748 3828 15804
rect 3828 15748 3832 15804
rect 3768 15744 3832 15748
rect 8680 15804 8744 15808
rect 8680 15748 8684 15804
rect 8684 15748 8740 15804
rect 8740 15748 8744 15804
rect 8680 15744 8744 15748
rect 8760 15804 8824 15808
rect 8760 15748 8764 15804
rect 8764 15748 8820 15804
rect 8820 15748 8824 15804
rect 8760 15744 8824 15748
rect 8840 15804 8904 15808
rect 8840 15748 8844 15804
rect 8844 15748 8900 15804
rect 8900 15748 8904 15804
rect 8840 15744 8904 15748
rect 8920 15804 8984 15808
rect 8920 15748 8924 15804
rect 8924 15748 8980 15804
rect 8980 15748 8984 15804
rect 8920 15744 8984 15748
rect 13832 15804 13896 15808
rect 13832 15748 13836 15804
rect 13836 15748 13892 15804
rect 13892 15748 13896 15804
rect 13832 15744 13896 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 6104 15260 6168 15264
rect 6104 15204 6108 15260
rect 6108 15204 6164 15260
rect 6164 15204 6168 15260
rect 6104 15200 6168 15204
rect 6184 15260 6248 15264
rect 6184 15204 6188 15260
rect 6188 15204 6244 15260
rect 6244 15204 6248 15260
rect 6184 15200 6248 15204
rect 6264 15260 6328 15264
rect 6264 15204 6268 15260
rect 6268 15204 6324 15260
rect 6324 15204 6328 15260
rect 6264 15200 6328 15204
rect 6344 15260 6408 15264
rect 6344 15204 6348 15260
rect 6348 15204 6404 15260
rect 6404 15204 6408 15260
rect 6344 15200 6408 15204
rect 11256 15260 11320 15264
rect 11256 15204 11260 15260
rect 11260 15204 11316 15260
rect 11316 15204 11320 15260
rect 11256 15200 11320 15204
rect 11336 15260 11400 15264
rect 11336 15204 11340 15260
rect 11340 15204 11396 15260
rect 11396 15204 11400 15260
rect 11336 15200 11400 15204
rect 11416 15260 11480 15264
rect 11416 15204 11420 15260
rect 11420 15204 11476 15260
rect 11476 15204 11480 15260
rect 11416 15200 11480 15204
rect 11496 15260 11560 15264
rect 11496 15204 11500 15260
rect 11500 15204 11556 15260
rect 11556 15204 11560 15260
rect 11496 15200 11560 15204
rect 3528 14716 3592 14720
rect 3528 14660 3532 14716
rect 3532 14660 3588 14716
rect 3588 14660 3592 14716
rect 3528 14656 3592 14660
rect 3608 14716 3672 14720
rect 3608 14660 3612 14716
rect 3612 14660 3668 14716
rect 3668 14660 3672 14716
rect 3608 14656 3672 14660
rect 3688 14716 3752 14720
rect 3688 14660 3692 14716
rect 3692 14660 3748 14716
rect 3748 14660 3752 14716
rect 3688 14656 3752 14660
rect 3768 14716 3832 14720
rect 3768 14660 3772 14716
rect 3772 14660 3828 14716
rect 3828 14660 3832 14716
rect 3768 14656 3832 14660
rect 8680 14716 8744 14720
rect 8680 14660 8684 14716
rect 8684 14660 8740 14716
rect 8740 14660 8744 14716
rect 8680 14656 8744 14660
rect 8760 14716 8824 14720
rect 8760 14660 8764 14716
rect 8764 14660 8820 14716
rect 8820 14660 8824 14716
rect 8760 14656 8824 14660
rect 8840 14716 8904 14720
rect 8840 14660 8844 14716
rect 8844 14660 8900 14716
rect 8900 14660 8904 14716
rect 8840 14656 8904 14660
rect 8920 14716 8984 14720
rect 8920 14660 8924 14716
rect 8924 14660 8980 14716
rect 8980 14660 8984 14716
rect 8920 14656 8984 14660
rect 13832 14716 13896 14720
rect 13832 14660 13836 14716
rect 13836 14660 13892 14716
rect 13892 14660 13896 14716
rect 13832 14656 13896 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 6104 14172 6168 14176
rect 6104 14116 6108 14172
rect 6108 14116 6164 14172
rect 6164 14116 6168 14172
rect 6104 14112 6168 14116
rect 6184 14172 6248 14176
rect 6184 14116 6188 14172
rect 6188 14116 6244 14172
rect 6244 14116 6248 14172
rect 6184 14112 6248 14116
rect 6264 14172 6328 14176
rect 6264 14116 6268 14172
rect 6268 14116 6324 14172
rect 6324 14116 6328 14172
rect 6264 14112 6328 14116
rect 6344 14172 6408 14176
rect 6344 14116 6348 14172
rect 6348 14116 6404 14172
rect 6404 14116 6408 14172
rect 6344 14112 6408 14116
rect 11256 14172 11320 14176
rect 11256 14116 11260 14172
rect 11260 14116 11316 14172
rect 11316 14116 11320 14172
rect 11256 14112 11320 14116
rect 11336 14172 11400 14176
rect 11336 14116 11340 14172
rect 11340 14116 11396 14172
rect 11396 14116 11400 14172
rect 11336 14112 11400 14116
rect 11416 14172 11480 14176
rect 11416 14116 11420 14172
rect 11420 14116 11476 14172
rect 11476 14116 11480 14172
rect 11416 14112 11480 14116
rect 11496 14172 11560 14176
rect 11496 14116 11500 14172
rect 11500 14116 11556 14172
rect 11556 14116 11560 14172
rect 11496 14112 11560 14116
rect 3528 13628 3592 13632
rect 3528 13572 3532 13628
rect 3532 13572 3588 13628
rect 3588 13572 3592 13628
rect 3528 13568 3592 13572
rect 3608 13628 3672 13632
rect 3608 13572 3612 13628
rect 3612 13572 3668 13628
rect 3668 13572 3672 13628
rect 3608 13568 3672 13572
rect 3688 13628 3752 13632
rect 3688 13572 3692 13628
rect 3692 13572 3748 13628
rect 3748 13572 3752 13628
rect 3688 13568 3752 13572
rect 3768 13628 3832 13632
rect 3768 13572 3772 13628
rect 3772 13572 3828 13628
rect 3828 13572 3832 13628
rect 3768 13568 3832 13572
rect 8680 13628 8744 13632
rect 8680 13572 8684 13628
rect 8684 13572 8740 13628
rect 8740 13572 8744 13628
rect 8680 13568 8744 13572
rect 8760 13628 8824 13632
rect 8760 13572 8764 13628
rect 8764 13572 8820 13628
rect 8820 13572 8824 13628
rect 8760 13568 8824 13572
rect 8840 13628 8904 13632
rect 8840 13572 8844 13628
rect 8844 13572 8900 13628
rect 8900 13572 8904 13628
rect 8840 13568 8904 13572
rect 8920 13628 8984 13632
rect 8920 13572 8924 13628
rect 8924 13572 8980 13628
rect 8980 13572 8984 13628
rect 8920 13568 8984 13572
rect 13832 13628 13896 13632
rect 13832 13572 13836 13628
rect 13836 13572 13892 13628
rect 13892 13572 13896 13628
rect 13832 13568 13896 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 6104 13084 6168 13088
rect 6104 13028 6108 13084
rect 6108 13028 6164 13084
rect 6164 13028 6168 13084
rect 6104 13024 6168 13028
rect 6184 13084 6248 13088
rect 6184 13028 6188 13084
rect 6188 13028 6244 13084
rect 6244 13028 6248 13084
rect 6184 13024 6248 13028
rect 6264 13084 6328 13088
rect 6264 13028 6268 13084
rect 6268 13028 6324 13084
rect 6324 13028 6328 13084
rect 6264 13024 6328 13028
rect 6344 13084 6408 13088
rect 6344 13028 6348 13084
rect 6348 13028 6404 13084
rect 6404 13028 6408 13084
rect 6344 13024 6408 13028
rect 11256 13084 11320 13088
rect 11256 13028 11260 13084
rect 11260 13028 11316 13084
rect 11316 13028 11320 13084
rect 11256 13024 11320 13028
rect 11336 13084 11400 13088
rect 11336 13028 11340 13084
rect 11340 13028 11396 13084
rect 11396 13028 11400 13084
rect 11336 13024 11400 13028
rect 11416 13084 11480 13088
rect 11416 13028 11420 13084
rect 11420 13028 11476 13084
rect 11476 13028 11480 13084
rect 11416 13024 11480 13028
rect 11496 13084 11560 13088
rect 11496 13028 11500 13084
rect 11500 13028 11556 13084
rect 11556 13028 11560 13084
rect 11496 13024 11560 13028
rect 3528 12540 3592 12544
rect 3528 12484 3532 12540
rect 3532 12484 3588 12540
rect 3588 12484 3592 12540
rect 3528 12480 3592 12484
rect 3608 12540 3672 12544
rect 3608 12484 3612 12540
rect 3612 12484 3668 12540
rect 3668 12484 3672 12540
rect 3608 12480 3672 12484
rect 3688 12540 3752 12544
rect 3688 12484 3692 12540
rect 3692 12484 3748 12540
rect 3748 12484 3752 12540
rect 3688 12480 3752 12484
rect 3768 12540 3832 12544
rect 3768 12484 3772 12540
rect 3772 12484 3828 12540
rect 3828 12484 3832 12540
rect 3768 12480 3832 12484
rect 8680 12540 8744 12544
rect 8680 12484 8684 12540
rect 8684 12484 8740 12540
rect 8740 12484 8744 12540
rect 8680 12480 8744 12484
rect 8760 12540 8824 12544
rect 8760 12484 8764 12540
rect 8764 12484 8820 12540
rect 8820 12484 8824 12540
rect 8760 12480 8824 12484
rect 8840 12540 8904 12544
rect 8840 12484 8844 12540
rect 8844 12484 8900 12540
rect 8900 12484 8904 12540
rect 8840 12480 8904 12484
rect 8920 12540 8984 12544
rect 8920 12484 8924 12540
rect 8924 12484 8980 12540
rect 8980 12484 8984 12540
rect 8920 12480 8984 12484
rect 13832 12540 13896 12544
rect 13832 12484 13836 12540
rect 13836 12484 13892 12540
rect 13892 12484 13896 12540
rect 13832 12480 13896 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 6104 11996 6168 12000
rect 6104 11940 6108 11996
rect 6108 11940 6164 11996
rect 6164 11940 6168 11996
rect 6104 11936 6168 11940
rect 6184 11996 6248 12000
rect 6184 11940 6188 11996
rect 6188 11940 6244 11996
rect 6244 11940 6248 11996
rect 6184 11936 6248 11940
rect 6264 11996 6328 12000
rect 6264 11940 6268 11996
rect 6268 11940 6324 11996
rect 6324 11940 6328 11996
rect 6264 11936 6328 11940
rect 6344 11996 6408 12000
rect 6344 11940 6348 11996
rect 6348 11940 6404 11996
rect 6404 11940 6408 11996
rect 6344 11936 6408 11940
rect 11256 11996 11320 12000
rect 11256 11940 11260 11996
rect 11260 11940 11316 11996
rect 11316 11940 11320 11996
rect 11256 11936 11320 11940
rect 11336 11996 11400 12000
rect 11336 11940 11340 11996
rect 11340 11940 11396 11996
rect 11396 11940 11400 11996
rect 11336 11936 11400 11940
rect 11416 11996 11480 12000
rect 11416 11940 11420 11996
rect 11420 11940 11476 11996
rect 11476 11940 11480 11996
rect 11416 11936 11480 11940
rect 11496 11996 11560 12000
rect 11496 11940 11500 11996
rect 11500 11940 11556 11996
rect 11556 11940 11560 11996
rect 11496 11936 11560 11940
rect 3528 11452 3592 11456
rect 3528 11396 3532 11452
rect 3532 11396 3588 11452
rect 3588 11396 3592 11452
rect 3528 11392 3592 11396
rect 3608 11452 3672 11456
rect 3608 11396 3612 11452
rect 3612 11396 3668 11452
rect 3668 11396 3672 11452
rect 3608 11392 3672 11396
rect 3688 11452 3752 11456
rect 3688 11396 3692 11452
rect 3692 11396 3748 11452
rect 3748 11396 3752 11452
rect 3688 11392 3752 11396
rect 3768 11452 3832 11456
rect 3768 11396 3772 11452
rect 3772 11396 3828 11452
rect 3828 11396 3832 11452
rect 3768 11392 3832 11396
rect 8680 11452 8744 11456
rect 8680 11396 8684 11452
rect 8684 11396 8740 11452
rect 8740 11396 8744 11452
rect 8680 11392 8744 11396
rect 8760 11452 8824 11456
rect 8760 11396 8764 11452
rect 8764 11396 8820 11452
rect 8820 11396 8824 11452
rect 8760 11392 8824 11396
rect 8840 11452 8904 11456
rect 8840 11396 8844 11452
rect 8844 11396 8900 11452
rect 8900 11396 8904 11452
rect 8840 11392 8904 11396
rect 8920 11452 8984 11456
rect 8920 11396 8924 11452
rect 8924 11396 8980 11452
rect 8980 11396 8984 11452
rect 8920 11392 8984 11396
rect 13832 11452 13896 11456
rect 13832 11396 13836 11452
rect 13836 11396 13892 11452
rect 13892 11396 13896 11452
rect 13832 11392 13896 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 6104 10908 6168 10912
rect 6104 10852 6108 10908
rect 6108 10852 6164 10908
rect 6164 10852 6168 10908
rect 6104 10848 6168 10852
rect 6184 10908 6248 10912
rect 6184 10852 6188 10908
rect 6188 10852 6244 10908
rect 6244 10852 6248 10908
rect 6184 10848 6248 10852
rect 6264 10908 6328 10912
rect 6264 10852 6268 10908
rect 6268 10852 6324 10908
rect 6324 10852 6328 10908
rect 6264 10848 6328 10852
rect 6344 10908 6408 10912
rect 6344 10852 6348 10908
rect 6348 10852 6404 10908
rect 6404 10852 6408 10908
rect 6344 10848 6408 10852
rect 11256 10908 11320 10912
rect 11256 10852 11260 10908
rect 11260 10852 11316 10908
rect 11316 10852 11320 10908
rect 11256 10848 11320 10852
rect 11336 10908 11400 10912
rect 11336 10852 11340 10908
rect 11340 10852 11396 10908
rect 11396 10852 11400 10908
rect 11336 10848 11400 10852
rect 11416 10908 11480 10912
rect 11416 10852 11420 10908
rect 11420 10852 11476 10908
rect 11476 10852 11480 10908
rect 11416 10848 11480 10852
rect 11496 10908 11560 10912
rect 11496 10852 11500 10908
rect 11500 10852 11556 10908
rect 11556 10852 11560 10908
rect 11496 10848 11560 10852
rect 3528 10364 3592 10368
rect 3528 10308 3532 10364
rect 3532 10308 3588 10364
rect 3588 10308 3592 10364
rect 3528 10304 3592 10308
rect 3608 10364 3672 10368
rect 3608 10308 3612 10364
rect 3612 10308 3668 10364
rect 3668 10308 3672 10364
rect 3608 10304 3672 10308
rect 3688 10364 3752 10368
rect 3688 10308 3692 10364
rect 3692 10308 3748 10364
rect 3748 10308 3752 10364
rect 3688 10304 3752 10308
rect 3768 10364 3832 10368
rect 3768 10308 3772 10364
rect 3772 10308 3828 10364
rect 3828 10308 3832 10364
rect 3768 10304 3832 10308
rect 8680 10364 8744 10368
rect 8680 10308 8684 10364
rect 8684 10308 8740 10364
rect 8740 10308 8744 10364
rect 8680 10304 8744 10308
rect 8760 10364 8824 10368
rect 8760 10308 8764 10364
rect 8764 10308 8820 10364
rect 8820 10308 8824 10364
rect 8760 10304 8824 10308
rect 8840 10364 8904 10368
rect 8840 10308 8844 10364
rect 8844 10308 8900 10364
rect 8900 10308 8904 10364
rect 8840 10304 8904 10308
rect 8920 10364 8984 10368
rect 8920 10308 8924 10364
rect 8924 10308 8980 10364
rect 8980 10308 8984 10364
rect 8920 10304 8984 10308
rect 13832 10364 13896 10368
rect 13832 10308 13836 10364
rect 13836 10308 13892 10364
rect 13892 10308 13896 10364
rect 13832 10304 13896 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 6104 9820 6168 9824
rect 6104 9764 6108 9820
rect 6108 9764 6164 9820
rect 6164 9764 6168 9820
rect 6104 9760 6168 9764
rect 6184 9820 6248 9824
rect 6184 9764 6188 9820
rect 6188 9764 6244 9820
rect 6244 9764 6248 9820
rect 6184 9760 6248 9764
rect 6264 9820 6328 9824
rect 6264 9764 6268 9820
rect 6268 9764 6324 9820
rect 6324 9764 6328 9820
rect 6264 9760 6328 9764
rect 6344 9820 6408 9824
rect 6344 9764 6348 9820
rect 6348 9764 6404 9820
rect 6404 9764 6408 9820
rect 6344 9760 6408 9764
rect 11256 9820 11320 9824
rect 11256 9764 11260 9820
rect 11260 9764 11316 9820
rect 11316 9764 11320 9820
rect 11256 9760 11320 9764
rect 11336 9820 11400 9824
rect 11336 9764 11340 9820
rect 11340 9764 11396 9820
rect 11396 9764 11400 9820
rect 11336 9760 11400 9764
rect 11416 9820 11480 9824
rect 11416 9764 11420 9820
rect 11420 9764 11476 9820
rect 11476 9764 11480 9820
rect 11416 9760 11480 9764
rect 11496 9820 11560 9824
rect 11496 9764 11500 9820
rect 11500 9764 11556 9820
rect 11556 9764 11560 9820
rect 11496 9760 11560 9764
rect 3528 9276 3592 9280
rect 3528 9220 3532 9276
rect 3532 9220 3588 9276
rect 3588 9220 3592 9276
rect 3528 9216 3592 9220
rect 3608 9276 3672 9280
rect 3608 9220 3612 9276
rect 3612 9220 3668 9276
rect 3668 9220 3672 9276
rect 3608 9216 3672 9220
rect 3688 9276 3752 9280
rect 3688 9220 3692 9276
rect 3692 9220 3748 9276
rect 3748 9220 3752 9276
rect 3688 9216 3752 9220
rect 3768 9276 3832 9280
rect 3768 9220 3772 9276
rect 3772 9220 3828 9276
rect 3828 9220 3832 9276
rect 3768 9216 3832 9220
rect 8680 9276 8744 9280
rect 8680 9220 8684 9276
rect 8684 9220 8740 9276
rect 8740 9220 8744 9276
rect 8680 9216 8744 9220
rect 8760 9276 8824 9280
rect 8760 9220 8764 9276
rect 8764 9220 8820 9276
rect 8820 9220 8824 9276
rect 8760 9216 8824 9220
rect 8840 9276 8904 9280
rect 8840 9220 8844 9276
rect 8844 9220 8900 9276
rect 8900 9220 8904 9276
rect 8840 9216 8904 9220
rect 8920 9276 8984 9280
rect 8920 9220 8924 9276
rect 8924 9220 8980 9276
rect 8980 9220 8984 9276
rect 8920 9216 8984 9220
rect 13832 9276 13896 9280
rect 13832 9220 13836 9276
rect 13836 9220 13892 9276
rect 13892 9220 13896 9276
rect 13832 9216 13896 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 6104 8732 6168 8736
rect 6104 8676 6108 8732
rect 6108 8676 6164 8732
rect 6164 8676 6168 8732
rect 6104 8672 6168 8676
rect 6184 8732 6248 8736
rect 6184 8676 6188 8732
rect 6188 8676 6244 8732
rect 6244 8676 6248 8732
rect 6184 8672 6248 8676
rect 6264 8732 6328 8736
rect 6264 8676 6268 8732
rect 6268 8676 6324 8732
rect 6324 8676 6328 8732
rect 6264 8672 6328 8676
rect 6344 8732 6408 8736
rect 6344 8676 6348 8732
rect 6348 8676 6404 8732
rect 6404 8676 6408 8732
rect 6344 8672 6408 8676
rect 11256 8732 11320 8736
rect 11256 8676 11260 8732
rect 11260 8676 11316 8732
rect 11316 8676 11320 8732
rect 11256 8672 11320 8676
rect 11336 8732 11400 8736
rect 11336 8676 11340 8732
rect 11340 8676 11396 8732
rect 11396 8676 11400 8732
rect 11336 8672 11400 8676
rect 11416 8732 11480 8736
rect 11416 8676 11420 8732
rect 11420 8676 11476 8732
rect 11476 8676 11480 8732
rect 11416 8672 11480 8676
rect 11496 8732 11560 8736
rect 11496 8676 11500 8732
rect 11500 8676 11556 8732
rect 11556 8676 11560 8732
rect 11496 8672 11560 8676
rect 3528 8188 3592 8192
rect 3528 8132 3532 8188
rect 3532 8132 3588 8188
rect 3588 8132 3592 8188
rect 3528 8128 3592 8132
rect 3608 8188 3672 8192
rect 3608 8132 3612 8188
rect 3612 8132 3668 8188
rect 3668 8132 3672 8188
rect 3608 8128 3672 8132
rect 3688 8188 3752 8192
rect 3688 8132 3692 8188
rect 3692 8132 3748 8188
rect 3748 8132 3752 8188
rect 3688 8128 3752 8132
rect 3768 8188 3832 8192
rect 3768 8132 3772 8188
rect 3772 8132 3828 8188
rect 3828 8132 3832 8188
rect 3768 8128 3832 8132
rect 8680 8188 8744 8192
rect 8680 8132 8684 8188
rect 8684 8132 8740 8188
rect 8740 8132 8744 8188
rect 8680 8128 8744 8132
rect 8760 8188 8824 8192
rect 8760 8132 8764 8188
rect 8764 8132 8820 8188
rect 8820 8132 8824 8188
rect 8760 8128 8824 8132
rect 8840 8188 8904 8192
rect 8840 8132 8844 8188
rect 8844 8132 8900 8188
rect 8900 8132 8904 8188
rect 8840 8128 8904 8132
rect 8920 8188 8984 8192
rect 8920 8132 8924 8188
rect 8924 8132 8980 8188
rect 8980 8132 8984 8188
rect 8920 8128 8984 8132
rect 13832 8188 13896 8192
rect 13832 8132 13836 8188
rect 13836 8132 13892 8188
rect 13892 8132 13896 8188
rect 13832 8128 13896 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 6104 7644 6168 7648
rect 6104 7588 6108 7644
rect 6108 7588 6164 7644
rect 6164 7588 6168 7644
rect 6104 7584 6168 7588
rect 6184 7644 6248 7648
rect 6184 7588 6188 7644
rect 6188 7588 6244 7644
rect 6244 7588 6248 7644
rect 6184 7584 6248 7588
rect 6264 7644 6328 7648
rect 6264 7588 6268 7644
rect 6268 7588 6324 7644
rect 6324 7588 6328 7644
rect 6264 7584 6328 7588
rect 6344 7644 6408 7648
rect 6344 7588 6348 7644
rect 6348 7588 6404 7644
rect 6404 7588 6408 7644
rect 6344 7584 6408 7588
rect 11256 7644 11320 7648
rect 11256 7588 11260 7644
rect 11260 7588 11316 7644
rect 11316 7588 11320 7644
rect 11256 7584 11320 7588
rect 11336 7644 11400 7648
rect 11336 7588 11340 7644
rect 11340 7588 11396 7644
rect 11396 7588 11400 7644
rect 11336 7584 11400 7588
rect 11416 7644 11480 7648
rect 11416 7588 11420 7644
rect 11420 7588 11476 7644
rect 11476 7588 11480 7644
rect 11416 7584 11480 7588
rect 11496 7644 11560 7648
rect 11496 7588 11500 7644
rect 11500 7588 11556 7644
rect 11556 7588 11560 7644
rect 11496 7584 11560 7588
rect 3528 7100 3592 7104
rect 3528 7044 3532 7100
rect 3532 7044 3588 7100
rect 3588 7044 3592 7100
rect 3528 7040 3592 7044
rect 3608 7100 3672 7104
rect 3608 7044 3612 7100
rect 3612 7044 3668 7100
rect 3668 7044 3672 7100
rect 3608 7040 3672 7044
rect 3688 7100 3752 7104
rect 3688 7044 3692 7100
rect 3692 7044 3748 7100
rect 3748 7044 3752 7100
rect 3688 7040 3752 7044
rect 3768 7100 3832 7104
rect 3768 7044 3772 7100
rect 3772 7044 3828 7100
rect 3828 7044 3832 7100
rect 3768 7040 3832 7044
rect 8680 7100 8744 7104
rect 8680 7044 8684 7100
rect 8684 7044 8740 7100
rect 8740 7044 8744 7100
rect 8680 7040 8744 7044
rect 8760 7100 8824 7104
rect 8760 7044 8764 7100
rect 8764 7044 8820 7100
rect 8820 7044 8824 7100
rect 8760 7040 8824 7044
rect 8840 7100 8904 7104
rect 8840 7044 8844 7100
rect 8844 7044 8900 7100
rect 8900 7044 8904 7100
rect 8840 7040 8904 7044
rect 8920 7100 8984 7104
rect 8920 7044 8924 7100
rect 8924 7044 8980 7100
rect 8980 7044 8984 7100
rect 8920 7040 8984 7044
rect 13832 7100 13896 7104
rect 13832 7044 13836 7100
rect 13836 7044 13892 7100
rect 13892 7044 13896 7100
rect 13832 7040 13896 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 6104 6556 6168 6560
rect 6104 6500 6108 6556
rect 6108 6500 6164 6556
rect 6164 6500 6168 6556
rect 6104 6496 6168 6500
rect 6184 6556 6248 6560
rect 6184 6500 6188 6556
rect 6188 6500 6244 6556
rect 6244 6500 6248 6556
rect 6184 6496 6248 6500
rect 6264 6556 6328 6560
rect 6264 6500 6268 6556
rect 6268 6500 6324 6556
rect 6324 6500 6328 6556
rect 6264 6496 6328 6500
rect 6344 6556 6408 6560
rect 6344 6500 6348 6556
rect 6348 6500 6404 6556
rect 6404 6500 6408 6556
rect 6344 6496 6408 6500
rect 11256 6556 11320 6560
rect 11256 6500 11260 6556
rect 11260 6500 11316 6556
rect 11316 6500 11320 6556
rect 11256 6496 11320 6500
rect 11336 6556 11400 6560
rect 11336 6500 11340 6556
rect 11340 6500 11396 6556
rect 11396 6500 11400 6556
rect 11336 6496 11400 6500
rect 11416 6556 11480 6560
rect 11416 6500 11420 6556
rect 11420 6500 11476 6556
rect 11476 6500 11480 6556
rect 11416 6496 11480 6500
rect 11496 6556 11560 6560
rect 11496 6500 11500 6556
rect 11500 6500 11556 6556
rect 11556 6500 11560 6556
rect 11496 6496 11560 6500
rect 3528 6012 3592 6016
rect 3528 5956 3532 6012
rect 3532 5956 3588 6012
rect 3588 5956 3592 6012
rect 3528 5952 3592 5956
rect 3608 6012 3672 6016
rect 3608 5956 3612 6012
rect 3612 5956 3668 6012
rect 3668 5956 3672 6012
rect 3608 5952 3672 5956
rect 3688 6012 3752 6016
rect 3688 5956 3692 6012
rect 3692 5956 3748 6012
rect 3748 5956 3752 6012
rect 3688 5952 3752 5956
rect 3768 6012 3832 6016
rect 3768 5956 3772 6012
rect 3772 5956 3828 6012
rect 3828 5956 3832 6012
rect 3768 5952 3832 5956
rect 8680 6012 8744 6016
rect 8680 5956 8684 6012
rect 8684 5956 8740 6012
rect 8740 5956 8744 6012
rect 8680 5952 8744 5956
rect 8760 6012 8824 6016
rect 8760 5956 8764 6012
rect 8764 5956 8820 6012
rect 8820 5956 8824 6012
rect 8760 5952 8824 5956
rect 8840 6012 8904 6016
rect 8840 5956 8844 6012
rect 8844 5956 8900 6012
rect 8900 5956 8904 6012
rect 8840 5952 8904 5956
rect 8920 6012 8984 6016
rect 8920 5956 8924 6012
rect 8924 5956 8980 6012
rect 8980 5956 8984 6012
rect 8920 5952 8984 5956
rect 13832 6012 13896 6016
rect 13832 5956 13836 6012
rect 13836 5956 13892 6012
rect 13892 5956 13896 6012
rect 13832 5952 13896 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 6104 5468 6168 5472
rect 6104 5412 6108 5468
rect 6108 5412 6164 5468
rect 6164 5412 6168 5468
rect 6104 5408 6168 5412
rect 6184 5468 6248 5472
rect 6184 5412 6188 5468
rect 6188 5412 6244 5468
rect 6244 5412 6248 5468
rect 6184 5408 6248 5412
rect 6264 5468 6328 5472
rect 6264 5412 6268 5468
rect 6268 5412 6324 5468
rect 6324 5412 6328 5468
rect 6264 5408 6328 5412
rect 6344 5468 6408 5472
rect 6344 5412 6348 5468
rect 6348 5412 6404 5468
rect 6404 5412 6408 5468
rect 6344 5408 6408 5412
rect 11256 5468 11320 5472
rect 11256 5412 11260 5468
rect 11260 5412 11316 5468
rect 11316 5412 11320 5468
rect 11256 5408 11320 5412
rect 11336 5468 11400 5472
rect 11336 5412 11340 5468
rect 11340 5412 11396 5468
rect 11396 5412 11400 5468
rect 11336 5408 11400 5412
rect 11416 5468 11480 5472
rect 11416 5412 11420 5468
rect 11420 5412 11476 5468
rect 11476 5412 11480 5468
rect 11416 5408 11480 5412
rect 11496 5468 11560 5472
rect 11496 5412 11500 5468
rect 11500 5412 11556 5468
rect 11556 5412 11560 5468
rect 11496 5408 11560 5412
rect 3528 4924 3592 4928
rect 3528 4868 3532 4924
rect 3532 4868 3588 4924
rect 3588 4868 3592 4924
rect 3528 4864 3592 4868
rect 3608 4924 3672 4928
rect 3608 4868 3612 4924
rect 3612 4868 3668 4924
rect 3668 4868 3672 4924
rect 3608 4864 3672 4868
rect 3688 4924 3752 4928
rect 3688 4868 3692 4924
rect 3692 4868 3748 4924
rect 3748 4868 3752 4924
rect 3688 4864 3752 4868
rect 3768 4924 3832 4928
rect 3768 4868 3772 4924
rect 3772 4868 3828 4924
rect 3828 4868 3832 4924
rect 3768 4864 3832 4868
rect 8680 4924 8744 4928
rect 8680 4868 8684 4924
rect 8684 4868 8740 4924
rect 8740 4868 8744 4924
rect 8680 4864 8744 4868
rect 8760 4924 8824 4928
rect 8760 4868 8764 4924
rect 8764 4868 8820 4924
rect 8820 4868 8824 4924
rect 8760 4864 8824 4868
rect 8840 4924 8904 4928
rect 8840 4868 8844 4924
rect 8844 4868 8900 4924
rect 8900 4868 8904 4924
rect 8840 4864 8904 4868
rect 8920 4924 8984 4928
rect 8920 4868 8924 4924
rect 8924 4868 8980 4924
rect 8980 4868 8984 4924
rect 8920 4864 8984 4868
rect 13832 4924 13896 4928
rect 13832 4868 13836 4924
rect 13836 4868 13892 4924
rect 13892 4868 13896 4924
rect 13832 4864 13896 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 6104 4380 6168 4384
rect 6104 4324 6108 4380
rect 6108 4324 6164 4380
rect 6164 4324 6168 4380
rect 6104 4320 6168 4324
rect 6184 4380 6248 4384
rect 6184 4324 6188 4380
rect 6188 4324 6244 4380
rect 6244 4324 6248 4380
rect 6184 4320 6248 4324
rect 6264 4380 6328 4384
rect 6264 4324 6268 4380
rect 6268 4324 6324 4380
rect 6324 4324 6328 4380
rect 6264 4320 6328 4324
rect 6344 4380 6408 4384
rect 6344 4324 6348 4380
rect 6348 4324 6404 4380
rect 6404 4324 6408 4380
rect 6344 4320 6408 4324
rect 11256 4380 11320 4384
rect 11256 4324 11260 4380
rect 11260 4324 11316 4380
rect 11316 4324 11320 4380
rect 11256 4320 11320 4324
rect 11336 4380 11400 4384
rect 11336 4324 11340 4380
rect 11340 4324 11396 4380
rect 11396 4324 11400 4380
rect 11336 4320 11400 4324
rect 11416 4380 11480 4384
rect 11416 4324 11420 4380
rect 11420 4324 11476 4380
rect 11476 4324 11480 4380
rect 11416 4320 11480 4324
rect 11496 4380 11560 4384
rect 11496 4324 11500 4380
rect 11500 4324 11556 4380
rect 11556 4324 11560 4380
rect 11496 4320 11560 4324
rect 3528 3836 3592 3840
rect 3528 3780 3532 3836
rect 3532 3780 3588 3836
rect 3588 3780 3592 3836
rect 3528 3776 3592 3780
rect 3608 3836 3672 3840
rect 3608 3780 3612 3836
rect 3612 3780 3668 3836
rect 3668 3780 3672 3836
rect 3608 3776 3672 3780
rect 3688 3836 3752 3840
rect 3688 3780 3692 3836
rect 3692 3780 3748 3836
rect 3748 3780 3752 3836
rect 3688 3776 3752 3780
rect 3768 3836 3832 3840
rect 3768 3780 3772 3836
rect 3772 3780 3828 3836
rect 3828 3780 3832 3836
rect 3768 3776 3832 3780
rect 8680 3836 8744 3840
rect 8680 3780 8684 3836
rect 8684 3780 8740 3836
rect 8740 3780 8744 3836
rect 8680 3776 8744 3780
rect 8760 3836 8824 3840
rect 8760 3780 8764 3836
rect 8764 3780 8820 3836
rect 8820 3780 8824 3836
rect 8760 3776 8824 3780
rect 8840 3836 8904 3840
rect 8840 3780 8844 3836
rect 8844 3780 8900 3836
rect 8900 3780 8904 3836
rect 8840 3776 8904 3780
rect 8920 3836 8984 3840
rect 8920 3780 8924 3836
rect 8924 3780 8980 3836
rect 8980 3780 8984 3836
rect 8920 3776 8984 3780
rect 13832 3836 13896 3840
rect 13832 3780 13836 3836
rect 13836 3780 13892 3836
rect 13892 3780 13896 3836
rect 13832 3776 13896 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 6104 3292 6168 3296
rect 6104 3236 6108 3292
rect 6108 3236 6164 3292
rect 6164 3236 6168 3292
rect 6104 3232 6168 3236
rect 6184 3292 6248 3296
rect 6184 3236 6188 3292
rect 6188 3236 6244 3292
rect 6244 3236 6248 3292
rect 6184 3232 6248 3236
rect 6264 3292 6328 3296
rect 6264 3236 6268 3292
rect 6268 3236 6324 3292
rect 6324 3236 6328 3292
rect 6264 3232 6328 3236
rect 6344 3292 6408 3296
rect 6344 3236 6348 3292
rect 6348 3236 6404 3292
rect 6404 3236 6408 3292
rect 6344 3232 6408 3236
rect 11256 3292 11320 3296
rect 11256 3236 11260 3292
rect 11260 3236 11316 3292
rect 11316 3236 11320 3292
rect 11256 3232 11320 3236
rect 11336 3292 11400 3296
rect 11336 3236 11340 3292
rect 11340 3236 11396 3292
rect 11396 3236 11400 3292
rect 11336 3232 11400 3236
rect 11416 3292 11480 3296
rect 11416 3236 11420 3292
rect 11420 3236 11476 3292
rect 11476 3236 11480 3292
rect 11416 3232 11480 3236
rect 11496 3292 11560 3296
rect 11496 3236 11500 3292
rect 11500 3236 11556 3292
rect 11556 3236 11560 3292
rect 11496 3232 11560 3236
rect 3528 2748 3592 2752
rect 3528 2692 3532 2748
rect 3532 2692 3588 2748
rect 3588 2692 3592 2748
rect 3528 2688 3592 2692
rect 3608 2748 3672 2752
rect 3608 2692 3612 2748
rect 3612 2692 3668 2748
rect 3668 2692 3672 2748
rect 3608 2688 3672 2692
rect 3688 2748 3752 2752
rect 3688 2692 3692 2748
rect 3692 2692 3748 2748
rect 3748 2692 3752 2748
rect 3688 2688 3752 2692
rect 3768 2748 3832 2752
rect 3768 2692 3772 2748
rect 3772 2692 3828 2748
rect 3828 2692 3832 2748
rect 3768 2688 3832 2692
rect 8680 2748 8744 2752
rect 8680 2692 8684 2748
rect 8684 2692 8740 2748
rect 8740 2692 8744 2748
rect 8680 2688 8744 2692
rect 8760 2748 8824 2752
rect 8760 2692 8764 2748
rect 8764 2692 8820 2748
rect 8820 2692 8824 2748
rect 8760 2688 8824 2692
rect 8840 2748 8904 2752
rect 8840 2692 8844 2748
rect 8844 2692 8900 2748
rect 8900 2692 8904 2748
rect 8840 2688 8904 2692
rect 8920 2748 8984 2752
rect 8920 2692 8924 2748
rect 8924 2692 8980 2748
rect 8980 2692 8984 2748
rect 8920 2688 8984 2692
rect 13832 2748 13896 2752
rect 13832 2692 13836 2748
rect 13836 2692 13892 2748
rect 13892 2692 13896 2748
rect 13832 2688 13896 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 6104 2204 6168 2208
rect 6104 2148 6108 2204
rect 6108 2148 6164 2204
rect 6164 2148 6168 2204
rect 6104 2144 6168 2148
rect 6184 2204 6248 2208
rect 6184 2148 6188 2204
rect 6188 2148 6244 2204
rect 6244 2148 6248 2204
rect 6184 2144 6248 2148
rect 6264 2204 6328 2208
rect 6264 2148 6268 2204
rect 6268 2148 6324 2204
rect 6324 2148 6328 2204
rect 6264 2144 6328 2148
rect 6344 2204 6408 2208
rect 6344 2148 6348 2204
rect 6348 2148 6404 2204
rect 6404 2148 6408 2204
rect 6344 2144 6408 2148
rect 11256 2204 11320 2208
rect 11256 2148 11260 2204
rect 11260 2148 11316 2204
rect 11316 2148 11320 2204
rect 11256 2144 11320 2148
rect 11336 2204 11400 2208
rect 11336 2148 11340 2204
rect 11340 2148 11396 2204
rect 11396 2148 11400 2204
rect 11336 2144 11400 2148
rect 11416 2204 11480 2208
rect 11416 2148 11420 2204
rect 11420 2148 11476 2204
rect 11476 2148 11480 2204
rect 11416 2144 11480 2148
rect 11496 2204 11560 2208
rect 11496 2148 11500 2204
rect 11500 2148 11556 2204
rect 11556 2148 11560 2204
rect 11496 2144 11560 2148
<< metal4 >>
rect 3520 16896 3840 17456
rect 3520 16832 3528 16896
rect 3592 16832 3608 16896
rect 3672 16832 3688 16896
rect 3752 16832 3768 16896
rect 3832 16832 3840 16896
rect 3520 15808 3840 16832
rect 3520 15744 3528 15808
rect 3592 15744 3608 15808
rect 3672 15744 3688 15808
rect 3752 15744 3768 15808
rect 3832 15744 3840 15808
rect 3520 14939 3840 15744
rect 3520 14720 3562 14939
rect 3798 14720 3840 14939
rect 3520 14656 3528 14720
rect 3592 14656 3608 14703
rect 3672 14656 3688 14703
rect 3752 14656 3768 14703
rect 3832 14656 3840 14720
rect 3520 13632 3840 14656
rect 3520 13568 3528 13632
rect 3592 13568 3608 13632
rect 3672 13568 3688 13632
rect 3752 13568 3768 13632
rect 3832 13568 3840 13632
rect 3520 12544 3840 13568
rect 3520 12480 3528 12544
rect 3592 12480 3608 12544
rect 3672 12480 3688 12544
rect 3752 12480 3768 12544
rect 3832 12480 3840 12544
rect 3520 11456 3840 12480
rect 3520 11392 3528 11456
rect 3592 11392 3608 11456
rect 3672 11392 3688 11456
rect 3752 11392 3768 11456
rect 3832 11392 3840 11456
rect 3520 10368 3840 11392
rect 3520 10304 3528 10368
rect 3592 10304 3608 10368
rect 3672 10304 3688 10368
rect 3752 10304 3768 10368
rect 3832 10304 3840 10368
rect 3520 9862 3840 10304
rect 3520 9626 3562 9862
rect 3798 9626 3840 9862
rect 3520 9280 3840 9626
rect 3520 9216 3528 9280
rect 3592 9216 3608 9280
rect 3672 9216 3688 9280
rect 3752 9216 3768 9280
rect 3832 9216 3840 9280
rect 3520 8192 3840 9216
rect 3520 8128 3528 8192
rect 3592 8128 3608 8192
rect 3672 8128 3688 8192
rect 3752 8128 3768 8192
rect 3832 8128 3840 8192
rect 3520 7104 3840 8128
rect 3520 7040 3528 7104
rect 3592 7040 3608 7104
rect 3672 7040 3688 7104
rect 3752 7040 3768 7104
rect 3832 7040 3840 7104
rect 3520 6016 3840 7040
rect 3520 5952 3528 6016
rect 3592 5952 3608 6016
rect 3672 5952 3688 6016
rect 3752 5952 3768 6016
rect 3832 5952 3840 6016
rect 3520 4928 3840 5952
rect 3520 4864 3528 4928
rect 3592 4864 3608 4928
rect 3672 4864 3688 4928
rect 3752 4864 3768 4928
rect 3832 4864 3840 4928
rect 3520 4784 3840 4864
rect 3520 4548 3562 4784
rect 3798 4548 3840 4784
rect 3520 3840 3840 4548
rect 3520 3776 3528 3840
rect 3592 3776 3608 3840
rect 3672 3776 3688 3840
rect 3752 3776 3768 3840
rect 3832 3776 3840 3840
rect 3520 2752 3840 3776
rect 3520 2688 3528 2752
rect 3592 2688 3608 2752
rect 3672 2688 3688 2752
rect 3752 2688 3768 2752
rect 3832 2688 3840 2752
rect 3520 2128 3840 2688
rect 6096 17440 6416 17456
rect 6096 17376 6104 17440
rect 6168 17376 6184 17440
rect 6248 17376 6264 17440
rect 6328 17376 6344 17440
rect 6408 17376 6416 17440
rect 6096 16352 6416 17376
rect 6096 16288 6104 16352
rect 6168 16288 6184 16352
rect 6248 16288 6264 16352
rect 6328 16288 6344 16352
rect 6408 16288 6416 16352
rect 6096 15264 6416 16288
rect 6096 15200 6104 15264
rect 6168 15200 6184 15264
rect 6248 15200 6264 15264
rect 6328 15200 6344 15264
rect 6408 15200 6416 15264
rect 6096 14176 6416 15200
rect 6096 14112 6104 14176
rect 6168 14112 6184 14176
rect 6248 14112 6264 14176
rect 6328 14112 6344 14176
rect 6408 14112 6416 14176
rect 6096 13088 6416 14112
rect 6096 13024 6104 13088
rect 6168 13024 6184 13088
rect 6248 13024 6264 13088
rect 6328 13024 6344 13088
rect 6408 13024 6416 13088
rect 6096 12400 6416 13024
rect 6096 12164 6138 12400
rect 6374 12164 6416 12400
rect 6096 12000 6416 12164
rect 6096 11936 6104 12000
rect 6168 11936 6184 12000
rect 6248 11936 6264 12000
rect 6328 11936 6344 12000
rect 6408 11936 6416 12000
rect 6096 10912 6416 11936
rect 6096 10848 6104 10912
rect 6168 10848 6184 10912
rect 6248 10848 6264 10912
rect 6328 10848 6344 10912
rect 6408 10848 6416 10912
rect 6096 9824 6416 10848
rect 6096 9760 6104 9824
rect 6168 9760 6184 9824
rect 6248 9760 6264 9824
rect 6328 9760 6344 9824
rect 6408 9760 6416 9824
rect 6096 8736 6416 9760
rect 6096 8672 6104 8736
rect 6168 8672 6184 8736
rect 6248 8672 6264 8736
rect 6328 8672 6344 8736
rect 6408 8672 6416 8736
rect 6096 7648 6416 8672
rect 6096 7584 6104 7648
rect 6168 7584 6184 7648
rect 6248 7584 6264 7648
rect 6328 7584 6344 7648
rect 6408 7584 6416 7648
rect 6096 7323 6416 7584
rect 6096 7087 6138 7323
rect 6374 7087 6416 7323
rect 6096 6560 6416 7087
rect 6096 6496 6104 6560
rect 6168 6496 6184 6560
rect 6248 6496 6264 6560
rect 6328 6496 6344 6560
rect 6408 6496 6416 6560
rect 6096 5472 6416 6496
rect 6096 5408 6104 5472
rect 6168 5408 6184 5472
rect 6248 5408 6264 5472
rect 6328 5408 6344 5472
rect 6408 5408 6416 5472
rect 6096 4384 6416 5408
rect 6096 4320 6104 4384
rect 6168 4320 6184 4384
rect 6248 4320 6264 4384
rect 6328 4320 6344 4384
rect 6408 4320 6416 4384
rect 6096 3296 6416 4320
rect 6096 3232 6104 3296
rect 6168 3232 6184 3296
rect 6248 3232 6264 3296
rect 6328 3232 6344 3296
rect 6408 3232 6416 3296
rect 6096 2208 6416 3232
rect 6096 2144 6104 2208
rect 6168 2144 6184 2208
rect 6248 2144 6264 2208
rect 6328 2144 6344 2208
rect 6408 2144 6416 2208
rect 6096 2128 6416 2144
rect 8672 16896 8992 17456
rect 8672 16832 8680 16896
rect 8744 16832 8760 16896
rect 8824 16832 8840 16896
rect 8904 16832 8920 16896
rect 8984 16832 8992 16896
rect 8672 15808 8992 16832
rect 8672 15744 8680 15808
rect 8744 15744 8760 15808
rect 8824 15744 8840 15808
rect 8904 15744 8920 15808
rect 8984 15744 8992 15808
rect 8672 14939 8992 15744
rect 8672 14720 8714 14939
rect 8950 14720 8992 14939
rect 8672 14656 8680 14720
rect 8744 14656 8760 14703
rect 8824 14656 8840 14703
rect 8904 14656 8920 14703
rect 8984 14656 8992 14720
rect 8672 13632 8992 14656
rect 8672 13568 8680 13632
rect 8744 13568 8760 13632
rect 8824 13568 8840 13632
rect 8904 13568 8920 13632
rect 8984 13568 8992 13632
rect 8672 12544 8992 13568
rect 8672 12480 8680 12544
rect 8744 12480 8760 12544
rect 8824 12480 8840 12544
rect 8904 12480 8920 12544
rect 8984 12480 8992 12544
rect 8672 11456 8992 12480
rect 8672 11392 8680 11456
rect 8744 11392 8760 11456
rect 8824 11392 8840 11456
rect 8904 11392 8920 11456
rect 8984 11392 8992 11456
rect 8672 10368 8992 11392
rect 8672 10304 8680 10368
rect 8744 10304 8760 10368
rect 8824 10304 8840 10368
rect 8904 10304 8920 10368
rect 8984 10304 8992 10368
rect 8672 9862 8992 10304
rect 8672 9626 8714 9862
rect 8950 9626 8992 9862
rect 8672 9280 8992 9626
rect 8672 9216 8680 9280
rect 8744 9216 8760 9280
rect 8824 9216 8840 9280
rect 8904 9216 8920 9280
rect 8984 9216 8992 9280
rect 8672 8192 8992 9216
rect 8672 8128 8680 8192
rect 8744 8128 8760 8192
rect 8824 8128 8840 8192
rect 8904 8128 8920 8192
rect 8984 8128 8992 8192
rect 8672 7104 8992 8128
rect 8672 7040 8680 7104
rect 8744 7040 8760 7104
rect 8824 7040 8840 7104
rect 8904 7040 8920 7104
rect 8984 7040 8992 7104
rect 8672 6016 8992 7040
rect 8672 5952 8680 6016
rect 8744 5952 8760 6016
rect 8824 5952 8840 6016
rect 8904 5952 8920 6016
rect 8984 5952 8992 6016
rect 8672 4928 8992 5952
rect 8672 4864 8680 4928
rect 8744 4864 8760 4928
rect 8824 4864 8840 4928
rect 8904 4864 8920 4928
rect 8984 4864 8992 4928
rect 8672 4784 8992 4864
rect 8672 4548 8714 4784
rect 8950 4548 8992 4784
rect 8672 3840 8992 4548
rect 8672 3776 8680 3840
rect 8744 3776 8760 3840
rect 8824 3776 8840 3840
rect 8904 3776 8920 3840
rect 8984 3776 8992 3840
rect 8672 2752 8992 3776
rect 8672 2688 8680 2752
rect 8744 2688 8760 2752
rect 8824 2688 8840 2752
rect 8904 2688 8920 2752
rect 8984 2688 8992 2752
rect 8672 2128 8992 2688
rect 11248 17440 11568 17456
rect 11248 17376 11256 17440
rect 11320 17376 11336 17440
rect 11400 17376 11416 17440
rect 11480 17376 11496 17440
rect 11560 17376 11568 17440
rect 11248 16352 11568 17376
rect 11248 16288 11256 16352
rect 11320 16288 11336 16352
rect 11400 16288 11416 16352
rect 11480 16288 11496 16352
rect 11560 16288 11568 16352
rect 11248 15264 11568 16288
rect 11248 15200 11256 15264
rect 11320 15200 11336 15264
rect 11400 15200 11416 15264
rect 11480 15200 11496 15264
rect 11560 15200 11568 15264
rect 11248 14176 11568 15200
rect 11248 14112 11256 14176
rect 11320 14112 11336 14176
rect 11400 14112 11416 14176
rect 11480 14112 11496 14176
rect 11560 14112 11568 14176
rect 11248 13088 11568 14112
rect 11248 13024 11256 13088
rect 11320 13024 11336 13088
rect 11400 13024 11416 13088
rect 11480 13024 11496 13088
rect 11560 13024 11568 13088
rect 11248 12400 11568 13024
rect 11248 12164 11290 12400
rect 11526 12164 11568 12400
rect 11248 12000 11568 12164
rect 11248 11936 11256 12000
rect 11320 11936 11336 12000
rect 11400 11936 11416 12000
rect 11480 11936 11496 12000
rect 11560 11936 11568 12000
rect 11248 10912 11568 11936
rect 11248 10848 11256 10912
rect 11320 10848 11336 10912
rect 11400 10848 11416 10912
rect 11480 10848 11496 10912
rect 11560 10848 11568 10912
rect 11248 9824 11568 10848
rect 11248 9760 11256 9824
rect 11320 9760 11336 9824
rect 11400 9760 11416 9824
rect 11480 9760 11496 9824
rect 11560 9760 11568 9824
rect 11248 8736 11568 9760
rect 11248 8672 11256 8736
rect 11320 8672 11336 8736
rect 11400 8672 11416 8736
rect 11480 8672 11496 8736
rect 11560 8672 11568 8736
rect 11248 7648 11568 8672
rect 11248 7584 11256 7648
rect 11320 7584 11336 7648
rect 11400 7584 11416 7648
rect 11480 7584 11496 7648
rect 11560 7584 11568 7648
rect 11248 7323 11568 7584
rect 11248 7087 11290 7323
rect 11526 7087 11568 7323
rect 11248 6560 11568 7087
rect 11248 6496 11256 6560
rect 11320 6496 11336 6560
rect 11400 6496 11416 6560
rect 11480 6496 11496 6560
rect 11560 6496 11568 6560
rect 11248 5472 11568 6496
rect 11248 5408 11256 5472
rect 11320 5408 11336 5472
rect 11400 5408 11416 5472
rect 11480 5408 11496 5472
rect 11560 5408 11568 5472
rect 11248 4384 11568 5408
rect 11248 4320 11256 4384
rect 11320 4320 11336 4384
rect 11400 4320 11416 4384
rect 11480 4320 11496 4384
rect 11560 4320 11568 4384
rect 11248 3296 11568 4320
rect 11248 3232 11256 3296
rect 11320 3232 11336 3296
rect 11400 3232 11416 3296
rect 11480 3232 11496 3296
rect 11560 3232 11568 3296
rect 11248 2208 11568 3232
rect 11248 2144 11256 2208
rect 11320 2144 11336 2208
rect 11400 2144 11416 2208
rect 11480 2144 11496 2208
rect 11560 2144 11568 2208
rect 11248 2128 11568 2144
rect 13824 16896 14144 17456
rect 13824 16832 13832 16896
rect 13896 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14144 16896
rect 13824 15808 14144 16832
rect 13824 15744 13832 15808
rect 13896 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14144 15808
rect 13824 14939 14144 15744
rect 13824 14720 13866 14939
rect 14102 14720 14144 14939
rect 13824 14656 13832 14720
rect 13896 14656 13912 14703
rect 13976 14656 13992 14703
rect 14056 14656 14072 14703
rect 14136 14656 14144 14720
rect 13824 13632 14144 14656
rect 13824 13568 13832 13632
rect 13896 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14144 13632
rect 13824 12544 14144 13568
rect 13824 12480 13832 12544
rect 13896 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14144 12544
rect 13824 11456 14144 12480
rect 13824 11392 13832 11456
rect 13896 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14144 11456
rect 13824 10368 14144 11392
rect 13824 10304 13832 10368
rect 13896 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14144 10368
rect 13824 9862 14144 10304
rect 13824 9626 13866 9862
rect 14102 9626 14144 9862
rect 13824 9280 14144 9626
rect 13824 9216 13832 9280
rect 13896 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14144 9280
rect 13824 8192 14144 9216
rect 13824 8128 13832 8192
rect 13896 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14144 8192
rect 13824 7104 14144 8128
rect 13824 7040 13832 7104
rect 13896 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14144 7104
rect 13824 6016 14144 7040
rect 13824 5952 13832 6016
rect 13896 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14144 6016
rect 13824 4928 14144 5952
rect 13824 4864 13832 4928
rect 13896 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14144 4928
rect 13824 4784 14144 4864
rect 13824 4548 13866 4784
rect 14102 4548 14144 4784
rect 13824 3840 14144 4548
rect 13824 3776 13832 3840
rect 13896 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14144 3840
rect 13824 2752 14144 3776
rect 13824 2688 13832 2752
rect 13896 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14144 2752
rect 13824 2128 14144 2688
<< via4 >>
rect 3562 14720 3798 14939
rect 3562 14703 3592 14720
rect 3592 14703 3608 14720
rect 3608 14703 3672 14720
rect 3672 14703 3688 14720
rect 3688 14703 3752 14720
rect 3752 14703 3768 14720
rect 3768 14703 3798 14720
rect 3562 9626 3798 9862
rect 3562 4548 3798 4784
rect 6138 12164 6374 12400
rect 6138 7087 6374 7323
rect 8714 14720 8950 14939
rect 8714 14703 8744 14720
rect 8744 14703 8760 14720
rect 8760 14703 8824 14720
rect 8824 14703 8840 14720
rect 8840 14703 8904 14720
rect 8904 14703 8920 14720
rect 8920 14703 8950 14720
rect 8714 9626 8950 9862
rect 8714 4548 8950 4784
rect 11290 12164 11526 12400
rect 11290 7087 11526 7323
rect 13866 14720 14102 14939
rect 13866 14703 13896 14720
rect 13896 14703 13912 14720
rect 13912 14703 13976 14720
rect 13976 14703 13992 14720
rect 13992 14703 14056 14720
rect 14056 14703 14072 14720
rect 14072 14703 14102 14720
rect 13866 9626 14102 9862
rect 13866 4548 14102 4784
<< metal5 >>
rect 1104 14939 16560 14981
rect 1104 14703 3562 14939
rect 3798 14703 8714 14939
rect 8950 14703 13866 14939
rect 14102 14703 16560 14939
rect 1104 14661 16560 14703
rect 1104 12400 16560 12442
rect 1104 12164 6138 12400
rect 6374 12164 11290 12400
rect 11526 12164 16560 12400
rect 1104 12122 16560 12164
rect 1104 9862 16560 9904
rect 1104 9626 3562 9862
rect 3798 9626 8714 9862
rect 8950 9626 13866 9862
rect 14102 9626 16560 9862
rect 1104 9584 16560 9626
rect 1104 7323 16560 7365
rect 1104 7087 6138 7323
rect 6374 7087 11290 7323
rect 11526 7087 16560 7323
rect 1104 7045 16560 7087
rect 1104 4784 16560 4827
rect 1104 4548 3562 4784
rect 3798 4548 8714 4784
rect 8950 4548 13866 4784
rect 14102 4548 16560 4784
rect 1104 4506 16560 4548
use sky130_fd_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1631199322
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1631199322
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1631199322
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1631199322
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1631199322
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1631199322
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1631199322
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31
timestamp 1631199322
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_sclk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 5888 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1631199322
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1631199322
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1631199322
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1631199322
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1631199322
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1631199322
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_60
timestamp 1631199322
transform 1 0 6624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 6532 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1631199322
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1631199322
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _17_
timestamp 1631199322
transform 1 0 7544 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 6992 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1631199322
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_84
timestamp 1631199322
transform 1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1631199322
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_93
timestamp 1631199322
transform 1 0 9660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1631199322
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_sclk
timestamp 1631199322
transform 1 0 9200 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__o22a_1  _13_
timestamp 1631199322
transform 1 0 10396 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1631199322
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1631199322
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1631199322
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1631199322
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1631199322
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1631199322
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1631199322
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1631199322
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _29_
timestamp 1631199322
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_1_133
timestamp 1631199322
transform 1 0 13340 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_145
timestamp 1631199322
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1631199322
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1631199322
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1631199322
transform -1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1631199322
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_161
timestamp 1631199322
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1631199322
transform -1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1631199322
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1631199322
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_149
timestamp 1631199322
transform 1 0 14812 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1631199322
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1631199322
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1631199322
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1631199322
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1631199322
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1631199322
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1631199322
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1631199322
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1631199322
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_45
timestamp 1631199322
transform 1 0 5244 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _18_
timestamp 1631199322
transform 1 0 5336 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _24_
timestamp 1631199322
transform 1 0 6348 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1631199322
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1631199322
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1631199322
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _26_
timestamp 1631199322
transform -1 0 10764 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1631199322
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _27_
timestamp 1631199322
transform 1 0 11132 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1631199322
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1631199322
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1631199322
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1631199322
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1631199322
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1631199322
transform -1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1631199322
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1631199322
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1631199322
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1631199322
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1631199322
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1631199322
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1631199322
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1631199322
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _23_
timestamp 1631199322
transform 1 0 6348 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_3_77
timestamp 1631199322
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_85
timestamp 1631199322
transform 1 0 8924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_sclk
timestamp 1631199322
transform 1 0 9016 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1631199322
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1631199322
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _14_
timestamp 1631199322
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _21_
timestamp 1631199322
transform 1 0 12512 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_3_106
timestamp 1631199322
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_131
timestamp 1631199322
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_143
timestamp 1631199322
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1631199322
transform -1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_155
timestamp 1631199322
transform 1 0 15364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1631199322
transform 1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1631199322
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1631199322
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1631199322
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1631199322
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1631199322
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1631199322
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1631199322
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_59
timestamp 1631199322
transform 1 0 6532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_53
timestamp 1631199322
transform 1 0 5980 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _22_
timestamp 1631199322
transform 1 0 6624 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1631199322
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_92
timestamp 1631199322
transform 1 0 9568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1631199322
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1631199322
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_1  _16_
timestamp 1631199322
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _28_
timestamp 1631199322
transform 1 0 10488 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_4_122
timestamp 1631199322
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1631199322
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1631199322
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1631199322
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1631199322
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1631199322
transform -1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1631199322
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1631199322
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1631199322
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1631199322
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1631199322
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1631199322
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1631199322
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1631199322
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1631199322
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_77
timestamp 1631199322
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_69
timestamp 1631199322
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _12_
timestamp 1631199322
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _20_
timestamp 1631199322
transform 1 0 7544 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_95
timestamp 1631199322
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1631199322
transform 1 0 8832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1631199322
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1631199322
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1631199322
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1631199322
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1631199322
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1631199322
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1631199322
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_161
timestamp 1631199322
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1631199322
transform -1 0 16560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1631199322
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1631199322
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1631199322
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1631199322
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1631199322
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1631199322
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1631199322
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1631199322
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1631199322
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1631199322
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1631199322
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1631199322
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1631199322
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1631199322
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1631199322
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1631199322
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1631199322
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1631199322
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1631199322
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1631199322
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1631199322
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1631199322
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1631199322
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1631199322
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1631199322
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1631199322
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1631199322
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1631199322
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1631199322
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1631199322
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1631199322
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1631199322
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1631199322
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1631199322
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1631199322
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1631199322
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1631199322
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1631199322
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1631199322
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1631199322
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_161
timestamp 1631199322
transform 1 0 15916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1631199322
transform -1 0 16560 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1631199322
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1631199322
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1631199322
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1631199322
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1631199322
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1631199322
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1631199322
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1631199322
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1631199322
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1631199322
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1631199322
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1631199322
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1631199322
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1631199322
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1631199322
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1631199322
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1631199322
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1631199322
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1631199322
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1631199322
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1631199322
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1631199322
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1631199322
transform -1 0 16560 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1631199322
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1631199322
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1631199322
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1631199322
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1631199322
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1631199322
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1631199322
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1631199322
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1631199322
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1631199322
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1631199322
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1631199322
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1631199322
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1631199322
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1631199322
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1631199322
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1631199322
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1631199322
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1631199322
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_161
timestamp 1631199322
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1631199322
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1631199322
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1631199322
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1631199322
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1631199322
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1631199322
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1631199322
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1631199322
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1631199322
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1631199322
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1631199322
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1631199322
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1631199322
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1631199322
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1631199322
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1631199322
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1631199322
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1631199322
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1631199322
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1631199322
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1631199322
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1631199322
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1631199322
transform -1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1631199322
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1631199322
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1631199322
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1631199322
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1631199322
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1631199322
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1631199322
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1631199322
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1631199322
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1631199322
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1631199322
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1631199322
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1631199322
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1631199322
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1631199322
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1631199322
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1631199322
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1631199322
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1631199322
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_161
timestamp 1631199322
transform 1 0 15916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1631199322
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1631199322
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1631199322
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1631199322
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1631199322
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1631199322
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1631199322
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1631199322
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1631199322
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1631199322
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1631199322
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1631199322
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1631199322
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1631199322
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1631199322
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1631199322
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1631199322
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1631199322
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1631199322
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1631199322
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1631199322
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1631199322
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1631199322
transform -1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1631199322
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1631199322
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1631199322
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1631199322
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1631199322
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1631199322
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1631199322
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1631199322
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1631199322
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1631199322
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1631199322
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1631199322
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1631199322
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1631199322
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1631199322
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1631199322
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1631199322
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1631199322
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1631199322
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1631199322
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1631199322
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1631199322
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1631199322
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1631199322
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1631199322
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1631199322
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1631199322
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1631199322
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1631199322
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1631199322
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1631199322
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1631199322
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1631199322
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1631199322
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1631199322
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1631199322
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1631199322
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1631199322
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1631199322
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1631199322
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_161
timestamp 1631199322
transform 1 0 15916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1631199322
transform -1 0 16560 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1631199322
transform -1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1631199322
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1631199322
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1631199322
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1631199322
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1631199322
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1631199322
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1631199322
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1631199322
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1631199322
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1631199322
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1631199322
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1631199322
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1631199322
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1631199322
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1631199322
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1631199322
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1631199322
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1631199322
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1631199322
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_161
timestamp 1631199322
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1631199322
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1631199322
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1631199322
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1631199322
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1631199322
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1631199322
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1631199322
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1631199322
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1631199322
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1631199322
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1631199322
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1631199322
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1631199322
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1631199322
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1631199322
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1631199322
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1631199322
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1631199322
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1631199322
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1631199322
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1631199322
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1631199322
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1631199322
transform -1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1631199322
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1631199322
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1631199322
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1631199322
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1631199322
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1631199322
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1631199322
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1631199322
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1631199322
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1631199322
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1631199322
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1631199322
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1631199322
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1631199322
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1631199322
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1631199322
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1631199322
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1631199322
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1631199322
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_161
timestamp 1631199322
transform 1 0 15916 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1631199322
transform -1 0 16560 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1631199322
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1631199322
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1631199322
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1631199322
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1631199322
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1631199322
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1631199322
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1631199322
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1631199322
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1631199322
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1631199322
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1631199322
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1631199322
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1631199322
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1631199322
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1631199322
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1631199322
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1631199322
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1631199322
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1631199322
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1631199322
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1631199322
transform -1 0 16560 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1631199322
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1631199322
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1631199322
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1631199322
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1631199322
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1631199322
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1631199322
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1631199322
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1631199322
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1631199322
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1631199322
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1631199322
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1631199322
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1631199322
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1631199322
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1631199322
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1631199322
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1631199322
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1631199322
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1631199322
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1631199322
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1631199322
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1631199322
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1631199322
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1631199322
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1631199322
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1631199322
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1631199322
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1631199322
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1631199322
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1631199322
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1631199322
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1631199322
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1631199322
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1631199322
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1631199322
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1631199322
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1631199322
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1631199322
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1631199322
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_161
timestamp 1631199322
transform 1 0 15916 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1631199322
transform -1 0 16560 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1631199322
transform -1 0 16560 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1631199322
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1631199322
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1631199322
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1631199322
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1631199322
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1631199322
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1631199322
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1631199322
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1631199322
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1631199322
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1631199322
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1631199322
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1631199322
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1631199322
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1631199322
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1631199322
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1631199322
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1631199322
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1631199322
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_161
timestamp 1631199322
transform 1 0 15916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1631199322
transform -1 0 16560 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1631199322
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1631199322
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1631199322
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1631199322
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1631199322
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1631199322
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1631199322
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1631199322
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1631199322
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1631199322
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1631199322
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1631199322
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1631199322
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1631199322
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1631199322
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1631199322
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1631199322
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1631199322
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1631199322
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1631199322
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1631199322
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1631199322
transform -1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1631199322
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1631199322
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1631199322
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1631199322
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1631199322
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1631199322
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1631199322
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1631199322
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1631199322
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1631199322
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1631199322
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1631199322
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1631199322
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1631199322
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1631199322
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1631199322
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1631199322
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1631199322
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1631199322
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_161
timestamp 1631199322
transform 1 0 15916 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1631199322
transform -1 0 16560 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1631199322
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1631199322
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1631199322
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1631199322
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1631199322
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1631199322
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1631199322
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1631199322
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1631199322
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1631199322
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1631199322
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1631199322
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1631199322
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1631199322
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1631199322
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1631199322
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1631199322
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1631199322
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1631199322
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1631199322
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1631199322
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1631199322
transform -1 0 16560 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1631199322
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1631199322
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1631199322
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1631199322
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1631199322
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1631199322
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1631199322
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1631199322
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1631199322
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1631199322
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1631199322
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1631199322
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1631199322
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1631199322
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1631199322
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1631199322
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1631199322
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1631199322
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1631199322
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_161
timestamp 1631199322
transform 1 0 15916 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1631199322
transform -1 0 16560 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1631199322
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1631199322
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1631199322
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1631199322
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1631199322
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_17
timestamp 1631199322
transform 1 0 2668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1631199322
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1631199322
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1631199322
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1631199322
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_29
timestamp 1631199322
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_41
timestamp 1631199322
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_25
timestamp 1631199322
transform 1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1631199322
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1631199322
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1631199322
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1631199322
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1631199322
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1631199322
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1631199322
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1631199322
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1631199322
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1631199322
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1631199322
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1631199322
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1631199322
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1631199322
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_85
timestamp 1631199322
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_97
timestamp 1631199322
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1631199322
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1631199322
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1631199322
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1631199322
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_116
timestamp 1631199322
transform 1 0 11776 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1631199322
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1631199322
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1631199322
transform -1 0 11776 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1631199322
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_128
timestamp 1631199322
transform 1 0 12880 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_141
timestamp 1631199322
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1631199322
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1631199322
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1631199322
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1631199322
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1631199322
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_161
timestamp 1631199322
transform 1 0 15916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1631199322
transform -1 0 16560 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1631199322
transform -1 0 16560 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1631199322
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 15364 0 -1 17408
box -38 -48 590 592
<< labels >>
rlabel metal5 s 1104 7045 16560 7365 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4507 16560 4827 6 VPWR
port 1 nsew power input
rlabel metal2 s 1122 0 1178 800 6 data[0]
port 2 nsew signal tristate
rlabel metal2 s 3330 0 3386 800 6 data[1]
port 3 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 data[2]
port 4 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 data[3]
port 5 nsew signal tristate
rlabel metal2 s 9954 0 10010 800 6 data[4]
port 6 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 data[5]
port 7 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 data[6]
port 8 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 data[7]
port 9 nsew signal tristate
rlabel metal2 s 15474 19084 15530 19884 6 reset
port 10 nsew signal input
rlabel metal2 s 6642 19084 6698 19884 6 sclk
port 11 nsew signal input
rlabel metal2 s 11058 19084 11114 19884 6 sdi
port 12 nsew signal input
rlabel metal2 s 2226 19084 2282 19884 6 ss
port 13 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 17740 19884
<< end >>
