magic
tech sky130A
magscale 1 2
timestamp 1634754066
<< metal1 >>
rect 3600 31840 3840 31980
rect 3600 31700 3660 31840
rect 3780 31700 3840 31840
rect 5840 31940 6100 31980
rect 5840 31800 5880 31940
rect 6000 31800 6100 31940
rect 5840 31760 6100 31800
rect 8300 31940 8520 31980
rect 8300 31800 8340 31940
rect 8460 31800 8520 31940
rect 8300 31740 8520 31800
rect 10580 31940 10880 31980
rect 10580 31800 10640 31940
rect 10760 31800 10880 31940
rect 10580 31700 10880 31800
rect 12880 31940 13120 31980
rect 12880 31800 12940 31940
rect 13060 31800 13120 31940
rect 12880 31760 13120 31800
rect 15220 31900 15460 31960
rect 15220 31760 15260 31900
rect 15380 31760 15460 31900
rect 15220 31720 15460 31760
rect 3600 31620 3840 31700
rect 10340 13480 10600 13660
rect 8540 13380 10600 13480
rect 6960 13180 7780 13380
rect 8020 13180 10600 13380
rect 8540 13080 10600 13180
rect 10340 12860 10600 13080
rect 10360 12840 10600 12860
rect 11900 12840 12240 13660
rect 13660 13280 13900 13640
rect 15020 13460 21620 13820
rect 13660 12920 17800 13280
rect 17520 12260 17800 12920
rect 17520 11900 21680 12260
rect 17520 10340 17800 11900
<< via1 >>
rect -900 31740 -780 31880
rect 1400 31760 1520 31900
rect 3660 31700 3780 31840
rect 5880 31800 6000 31940
rect 8340 31800 8460 31940
rect 10640 31800 10760 31940
rect 12940 31800 13060 31940
rect 15260 31760 15380 31900
<< metal2 >>
rect -940 31880 -740 35620
rect -940 31740 -900 31880
rect -780 31740 -740 31880
rect -940 31700 -740 31740
rect 1360 31900 1560 35640
rect 1360 31760 1400 31900
rect 1520 31760 1560 31900
rect 1360 31720 1560 31760
rect 3600 31840 3820 35600
rect 3600 31700 3660 31840
rect 3780 31700 3820 31840
rect 5840 31940 6040 35680
rect 5840 31800 5880 31940
rect 6000 31800 6040 31940
rect 5840 31760 6040 31800
rect 8300 31940 8500 35700
rect 8300 31800 8340 31940
rect 8460 31800 8500 31940
rect 8300 31740 8500 31800
rect 10600 31940 10800 35680
rect 10600 31800 10640 31940
rect 10760 31800 10800 31940
rect 10600 31760 10800 31800
rect 12900 31940 13100 35680
rect 15240 31960 15440 35660
rect 12900 31800 12940 31940
rect 13060 31800 13100 31940
rect 12900 31760 13100 31800
rect 15220 31900 15460 31960
rect 15220 31760 15260 31900
rect 15380 31760 15460 31900
rect 15220 31720 15460 31760
rect 3600 31620 3820 31700
use sky130_fd_pr__res_high_po_0p35_LN2BL5  XRI
timestamp 1634754066
transform 0 -1 7906 1 0 13275
box -201 -696 201 696
use digpot  digpot_0 ~/sky130_skel/dpga-ieee-sscs-contest-main/magic/digpot/mag
timestamp 1634754066
transform 1 0 1172 0 1 -1182
box -2100 14620 15416 33360
use ota  ota_0 ~/sky130_skel/dpga-ieee-sscs-contest-main/magic/ota/mag
timestamp 1634750299
transform 1 0 10840 0 1 3200
box -1120 -300 6960 9860
use spi_slave  spi_slave_0 ~/sky130_skel/dpga-ieee-sscs-contest-main/magic/spi/magic
timestamp 1634602588
transform 1 0 -2046 0 1 34420
box 1066 0 17518 20731
<< end >>
