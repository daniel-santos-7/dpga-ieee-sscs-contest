magic
tech sky130A
timestamp 1622553964
<< nwell >>
rect 4955 1385 5080 1735
rect 5210 1235 5335 1585
rect 5700 1385 5825 1735
rect 5955 1235 6080 1585
rect 6305 1385 6430 1735
rect 6970 1715 7110 1830
rect 7565 1715 7705 1830
rect 6560 1235 6685 1585
rect 6970 1550 7095 1715
rect 7225 1550 7350 1590
rect 6970 1390 7350 1550
rect 7565 1550 7690 1715
rect 7820 1550 7945 1590
rect 7565 1390 7945 1550
rect 7225 1240 7350 1390
rect 7820 1240 7945 1390
rect 4950 940 5090 1055
rect 5695 940 5835 1055
rect 6300 940 6440 1055
rect 6965 945 7105 1060
rect 7560 945 7700 1060
rect 4950 775 5075 940
rect 5205 775 5330 815
rect 4950 615 5330 775
rect 5695 775 5820 940
rect 5950 775 6075 815
rect 5695 615 6075 775
rect 6300 775 6425 940
rect 6555 775 6680 815
rect 6300 615 6680 775
rect 6965 780 7090 945
rect 7220 780 7345 820
rect 6965 620 7345 780
rect 7560 780 7685 945
rect 9170 890 10920 1790
rect 7815 780 7940 820
rect 7560 620 7940 780
rect 5205 465 5330 615
rect 5950 465 6075 615
rect 6555 465 6680 615
rect 7220 470 7345 620
rect 7815 470 7940 620
rect 9170 330 9920 890
rect 10570 651 10920 890
rect 4950 -195 5075 155
rect 5205 -345 5330 5
rect 5695 -195 5820 155
rect 5950 -345 6075 5
rect 6300 -195 6425 155
rect 6555 -345 6680 5
rect 6965 -190 7090 160
rect 7560 135 7700 250
rect 7220 -340 7345 10
rect 7560 -30 7685 135
rect 10570 21 11070 651
rect 7815 -30 7940 10
rect 7560 -190 7940 -30
rect 7815 -340 7940 -190
<< nmos >>
rect 5265 1620 5280 1720
rect 5010 1235 5025 1335
rect 5260 850 5275 950
rect 5005 465 5020 565
rect 5260 40 5275 140
rect 6010 1620 6025 1720
rect 5755 1235 5770 1335
rect 6615 1620 6630 1720
rect 6005 850 6020 950
rect 5750 465 5765 565
rect 6360 1235 6375 1335
rect 7280 1625 7295 1725
rect 6610 850 6625 950
rect 7025 1240 7040 1340
rect 7875 1625 7890 1725
rect 7620 1240 7635 1340
rect 6355 465 6370 565
rect 7275 855 7290 955
rect 7020 470 7035 570
rect 7870 855 7885 955
rect 5005 -345 5020 -245
rect 6005 40 6020 140
rect 7615 470 7630 570
rect 5750 -345 5765 -245
rect 6610 40 6625 140
rect 6355 -345 6370 -245
rect 7275 45 7290 145
rect 7020 -340 7035 -240
rect 7870 45 7885 145
rect 7615 -340 7630 -240
rect 9270 -70 9370 16
rect 9420 -70 9520 16
rect 9570 -70 9670 16
rect 9720 -70 9820 16
rect 10040 -210 10140 651
rect 10190 -210 10290 651
rect 10340 -210 10440 651
<< pmos >>
rect 5010 1410 5025 1710
rect 5265 1260 5280 1560
rect 5005 640 5020 940
rect 5260 490 5275 790
rect 5005 -170 5020 130
rect 5755 1410 5770 1710
rect 6010 1260 6025 1560
rect 6360 1410 6375 1710
rect 5750 640 5765 940
rect 6005 490 6020 790
rect 6615 1260 6630 1560
rect 7025 1415 7040 1715
rect 6355 640 6370 940
rect 7280 1265 7295 1565
rect 7620 1415 7635 1715
rect 7875 1265 7890 1565
rect 6610 490 6625 790
rect 7020 645 7035 945
rect 7275 495 7290 795
rect 7615 645 7630 945
rect 9270 940 9370 1525
rect 9420 940 9520 1525
rect 9570 940 9670 1525
rect 9820 940 9920 1525
rect 9970 940 10070 1525
rect 10120 940 10220 1525
rect 10270 940 10370 1525
rect 10420 940 10520 1525
rect 10570 940 10670 1525
rect 10720 940 10820 1525
rect 5260 -320 5275 -20
rect 5750 -170 5765 130
rect 7870 495 7885 795
rect 9270 380 9370 673
rect 9420 380 9520 673
rect 9570 380 9670 673
rect 9720 380 9820 673
rect 6005 -320 6020 -20
rect 6355 -170 6370 130
rect 6610 -320 6625 -20
rect 7020 -165 7035 135
rect 7275 -315 7290 -15
rect 7615 -165 7630 135
rect 7870 -315 7885 -15
rect 10620 41 10720 626
rect 10770 41 10870 626
rect 10920 41 11020 626
<< ndiff >>
rect 5230 1620 5265 1720
rect 5280 1620 5315 1720
rect 4975 1235 5010 1335
rect 5025 1235 5060 1335
rect 5225 940 5260 950
rect 5225 910 5230 940
rect 5250 910 5260 940
rect 5225 890 5260 910
rect 5225 860 5230 890
rect 5250 860 5260 890
rect 5225 850 5260 860
rect 5275 940 5310 950
rect 5275 910 5285 940
rect 5305 910 5310 940
rect 5275 890 5310 910
rect 5275 860 5285 890
rect 5305 860 5310 890
rect 5275 850 5310 860
rect 4970 555 5005 565
rect 4970 525 4975 555
rect 4995 525 5005 555
rect 4970 505 5005 525
rect 4970 475 4975 505
rect 4995 475 5005 505
rect 4970 465 5005 475
rect 5020 555 5055 565
rect 5020 525 5030 555
rect 5050 525 5055 555
rect 5020 505 5055 525
rect 5020 475 5030 505
rect 5050 475 5055 505
rect 5020 465 5055 475
rect 5225 40 5260 140
rect 5275 40 5310 140
rect 5975 1620 6010 1720
rect 6025 1620 6060 1720
rect 5720 1235 5755 1335
rect 5770 1235 5805 1335
rect 6580 1620 6615 1720
rect 6630 1620 6665 1720
rect 7245 1715 7280 1725
rect 5970 940 6005 950
rect 5970 910 5975 940
rect 5995 910 6005 940
rect 5970 890 6005 910
rect 5970 860 5975 890
rect 5995 860 6005 890
rect 5970 850 6005 860
rect 6020 940 6055 950
rect 6020 910 6030 940
rect 6050 910 6055 940
rect 6020 890 6055 910
rect 6020 860 6030 890
rect 6050 860 6055 890
rect 6020 850 6055 860
rect 5715 555 5750 565
rect 5715 525 5720 555
rect 5740 525 5750 555
rect 5715 505 5750 525
rect 5715 475 5720 505
rect 5740 475 5750 505
rect 5715 465 5750 475
rect 5765 555 5800 565
rect 5765 525 5775 555
rect 5795 525 5800 555
rect 5765 505 5800 525
rect 5765 475 5775 505
rect 5795 475 5800 505
rect 5765 465 5800 475
rect 6325 1235 6360 1335
rect 6375 1235 6410 1335
rect 7245 1685 7250 1715
rect 7270 1685 7280 1715
rect 7245 1665 7280 1685
rect 7245 1635 7250 1665
rect 7270 1635 7280 1665
rect 7245 1625 7280 1635
rect 7295 1715 7330 1725
rect 7840 1715 7875 1725
rect 7295 1685 7305 1715
rect 7325 1685 7330 1715
rect 7295 1665 7330 1685
rect 7295 1635 7305 1665
rect 7325 1635 7330 1665
rect 7295 1625 7330 1635
rect 6575 940 6610 950
rect 6575 910 6580 940
rect 6600 910 6610 940
rect 6575 890 6610 910
rect 6575 860 6580 890
rect 6600 860 6610 890
rect 6575 850 6610 860
rect 6625 940 6660 950
rect 6625 910 6635 940
rect 6655 910 6660 940
rect 6625 890 6660 910
rect 6625 860 6635 890
rect 6655 860 6660 890
rect 6625 850 6660 860
rect 6990 1330 7025 1340
rect 6990 1300 6995 1330
rect 7015 1300 7025 1330
rect 6990 1280 7025 1300
rect 6990 1250 6995 1280
rect 7015 1250 7025 1280
rect 6990 1240 7025 1250
rect 7040 1330 7075 1340
rect 7040 1300 7050 1330
rect 7070 1300 7075 1330
rect 7040 1280 7075 1300
rect 7040 1250 7050 1280
rect 7070 1250 7075 1280
rect 7840 1685 7845 1715
rect 7865 1685 7875 1715
rect 7840 1665 7875 1685
rect 7840 1635 7845 1665
rect 7865 1635 7875 1665
rect 7840 1625 7875 1635
rect 7890 1715 7925 1725
rect 7890 1685 7900 1715
rect 7920 1685 7925 1715
rect 7890 1665 7925 1685
rect 7890 1635 7900 1665
rect 7920 1635 7925 1665
rect 7890 1625 7925 1635
rect 7040 1240 7075 1250
rect 7585 1330 7620 1340
rect 7585 1300 7590 1330
rect 7610 1300 7620 1330
rect 7585 1280 7620 1300
rect 7585 1250 7590 1280
rect 7610 1250 7620 1280
rect 7585 1240 7620 1250
rect 7635 1330 7670 1340
rect 7635 1300 7645 1330
rect 7665 1300 7670 1330
rect 7635 1280 7670 1300
rect 7635 1250 7645 1280
rect 7665 1250 7670 1280
rect 7635 1240 7670 1250
rect 7240 945 7275 955
rect 6320 555 6355 565
rect 6320 525 6325 555
rect 6345 525 6355 555
rect 6320 505 6355 525
rect 6320 475 6325 505
rect 6345 475 6355 505
rect 6320 465 6355 475
rect 6370 555 6405 565
rect 6370 525 6380 555
rect 6400 525 6405 555
rect 6370 505 6405 525
rect 6370 475 6380 505
rect 6400 475 6405 505
rect 7240 915 7245 945
rect 7265 915 7275 945
rect 7240 895 7275 915
rect 7240 865 7245 895
rect 7265 865 7275 895
rect 7240 855 7275 865
rect 7290 945 7325 955
rect 7835 945 7870 955
rect 7290 915 7300 945
rect 7320 915 7325 945
rect 7290 895 7325 915
rect 7290 865 7300 895
rect 7320 865 7325 895
rect 7290 855 7325 865
rect 6985 560 7020 570
rect 6985 530 6990 560
rect 7010 530 7020 560
rect 6985 510 7020 530
rect 6370 465 6405 475
rect 6985 480 6990 510
rect 7010 480 7020 510
rect 6985 470 7020 480
rect 7035 560 7070 570
rect 7035 530 7045 560
rect 7065 530 7070 560
rect 7035 510 7070 530
rect 7035 480 7045 510
rect 7065 480 7070 510
rect 7835 915 7840 945
rect 7860 915 7870 945
rect 7835 895 7870 915
rect 7835 865 7840 895
rect 7860 865 7870 895
rect 7835 855 7870 865
rect 7885 945 7920 955
rect 7885 915 7895 945
rect 7915 915 7920 945
rect 7885 895 7920 915
rect 7885 865 7895 895
rect 7915 865 7920 895
rect 7885 855 7920 865
rect 7035 470 7070 480
rect 4970 -345 5005 -245
rect 5020 -345 5055 -245
rect 5970 40 6005 140
rect 6020 40 6055 140
rect 7580 560 7615 570
rect 7580 530 7585 560
rect 7605 530 7615 560
rect 7580 510 7615 530
rect 7580 480 7585 510
rect 7605 480 7615 510
rect 7580 470 7615 480
rect 7630 560 7665 570
rect 7630 530 7640 560
rect 7660 530 7665 560
rect 7630 510 7665 530
rect 7630 480 7640 510
rect 7660 480 7665 510
rect 7630 470 7665 480
rect 5715 -345 5750 -245
rect 5765 -345 5800 -245
rect 6575 40 6610 140
rect 6625 40 6660 140
rect 6320 -345 6355 -245
rect 6370 -345 6405 -245
rect 7240 45 7275 145
rect 7290 45 7325 145
rect 7835 135 7870 145
rect 6985 -340 7020 -240
rect 7035 -340 7070 -240
rect 7835 105 7840 135
rect 7860 105 7870 135
rect 7835 85 7870 105
rect 7835 55 7840 85
rect 7860 55 7870 85
rect 7835 45 7870 55
rect 7885 135 7920 145
rect 7885 105 7895 135
rect 7915 105 7920 135
rect 7885 85 7920 105
rect 7885 55 7895 85
rect 7915 55 7920 85
rect 7885 45 7920 55
rect 7580 -250 7615 -240
rect 7580 -280 7585 -250
rect 7605 -280 7615 -250
rect 7580 -300 7615 -280
rect 7580 -330 7585 -300
rect 7605 -330 7615 -300
rect 7580 -340 7615 -330
rect 7630 -250 7665 -240
rect 7630 -280 7640 -250
rect 7660 -280 7665 -250
rect 7630 -300 7665 -280
rect 7630 -330 7640 -300
rect 7660 -330 7665 -300
rect 9220 -70 9270 16
rect 9370 0 9420 16
rect 9370 -50 9380 0
rect 9410 -50 9420 0
rect 9370 -70 9420 -50
rect 9520 0 9570 16
rect 9520 -50 9530 0
rect 9560 -50 9570 0
rect 9520 -70 9570 -50
rect 9670 0 9720 16
rect 9670 -50 9680 0
rect 9710 -50 9720 0
rect 9670 -70 9720 -50
rect 9820 -70 9870 16
rect 9990 -210 10040 651
rect 10140 630 10190 651
rect 10140 600 10150 630
rect 10180 600 10190 630
rect 10140 580 10190 600
rect 10140 550 10150 580
rect 10180 550 10190 580
rect 10140 530 10190 550
rect 10140 500 10150 530
rect 10180 500 10190 530
rect 10140 480 10190 500
rect 10140 450 10150 480
rect 10180 450 10190 480
rect 10140 430 10190 450
rect 10140 400 10150 430
rect 10180 400 10190 430
rect 10140 380 10190 400
rect 10140 350 10150 380
rect 10180 350 10190 380
rect 10140 330 10190 350
rect 10140 300 10150 330
rect 10180 300 10190 330
rect 10140 280 10190 300
rect 10140 250 10150 280
rect 10180 250 10190 280
rect 10140 230 10190 250
rect 10140 200 10150 230
rect 10180 200 10190 230
rect 10140 180 10190 200
rect 10140 150 10150 180
rect 10180 150 10190 180
rect 10140 130 10190 150
rect 10140 100 10150 130
rect 10180 100 10190 130
rect 10140 80 10190 100
rect 10140 50 10150 80
rect 10180 50 10190 80
rect 10140 30 10190 50
rect 10140 0 10150 30
rect 10180 0 10190 30
rect 10140 -20 10190 0
rect 10140 -50 10150 -20
rect 10180 -50 10190 -20
rect 10140 -70 10190 -50
rect 10140 -100 10150 -70
rect 10180 -100 10190 -70
rect 10140 -120 10190 -100
rect 10140 -150 10150 -120
rect 10180 -150 10190 -120
rect 10140 -170 10190 -150
rect 10140 -200 10150 -170
rect 10180 -200 10190 -170
rect 10140 -210 10190 -200
rect 10290 630 10340 651
rect 10290 600 10300 630
rect 10330 600 10340 630
rect 10290 580 10340 600
rect 10290 550 10300 580
rect 10330 550 10340 580
rect 10290 530 10340 550
rect 10290 500 10300 530
rect 10330 500 10340 530
rect 10290 480 10340 500
rect 10290 450 10300 480
rect 10330 450 10340 480
rect 10290 430 10340 450
rect 10290 400 10300 430
rect 10330 400 10340 430
rect 10290 380 10340 400
rect 10290 350 10300 380
rect 10330 350 10340 380
rect 10290 330 10340 350
rect 10290 300 10300 330
rect 10330 300 10340 330
rect 10290 280 10340 300
rect 10290 250 10300 280
rect 10330 250 10340 280
rect 10290 230 10340 250
rect 10290 200 10300 230
rect 10330 200 10340 230
rect 10290 180 10340 200
rect 10290 150 10300 180
rect 10330 150 10340 180
rect 10290 130 10340 150
rect 10290 100 10300 130
rect 10330 100 10340 130
rect 10290 80 10340 100
rect 10290 50 10300 80
rect 10330 50 10340 80
rect 10290 30 10340 50
rect 10290 0 10300 30
rect 10330 0 10340 30
rect 10290 -20 10340 0
rect 10290 -50 10300 -20
rect 10330 -50 10340 -20
rect 10290 -70 10340 -50
rect 10290 -100 10300 -70
rect 10330 -100 10340 -70
rect 10290 -120 10340 -100
rect 10290 -150 10300 -120
rect 10330 -150 10340 -120
rect 10290 -170 10340 -150
rect 10290 -200 10300 -170
rect 10330 -200 10340 -170
rect 10290 -210 10340 -200
rect 10440 -210 10490 651
rect 7630 -340 7665 -330
<< pdiff >>
rect 4975 1410 5010 1710
rect 5025 1410 5060 1710
rect 5230 1260 5265 1560
rect 5280 1260 5315 1560
rect 4970 930 5005 940
rect 4970 900 4975 930
rect 4995 900 5005 930
rect 4970 865 5005 900
rect 4970 835 4975 865
rect 4995 835 5005 865
rect 4970 805 5005 835
rect 4970 775 4975 805
rect 4995 775 5005 805
rect 4970 740 5005 775
rect 4970 710 4975 740
rect 4995 710 5005 740
rect 4970 680 5005 710
rect 4970 650 4975 680
rect 4995 650 5005 680
rect 4970 640 5005 650
rect 5020 930 5055 940
rect 5020 900 5030 930
rect 5050 900 5055 930
rect 5020 870 5055 900
rect 5020 840 5030 870
rect 5050 840 5055 870
rect 5020 805 5055 840
rect 5020 775 5030 805
rect 5050 775 5055 805
rect 5020 745 5055 775
rect 5020 715 5030 745
rect 5050 715 5055 745
rect 5020 680 5055 715
rect 5020 650 5030 680
rect 5050 650 5055 680
rect 5020 640 5055 650
rect 5225 780 5260 790
rect 5225 750 5230 780
rect 5250 750 5260 780
rect 5225 715 5260 750
rect 5225 685 5230 715
rect 5250 685 5260 715
rect 5225 655 5260 685
rect 5225 625 5230 655
rect 5250 625 5260 655
rect 5225 590 5260 625
rect 5225 560 5230 590
rect 5250 560 5260 590
rect 5225 530 5260 560
rect 5225 500 5230 530
rect 5250 500 5260 530
rect 5225 490 5260 500
rect 5275 780 5310 790
rect 5275 750 5285 780
rect 5305 750 5310 780
rect 5275 720 5310 750
rect 5275 690 5285 720
rect 5305 690 5310 720
rect 5275 655 5310 690
rect 5275 625 5285 655
rect 5305 625 5310 655
rect 5275 595 5310 625
rect 5275 565 5285 595
rect 5305 565 5310 595
rect 5275 530 5310 565
rect 5275 500 5285 530
rect 5305 500 5310 530
rect 5275 490 5310 500
rect 4970 -170 5005 130
rect 5020 -170 5055 130
rect 5720 1410 5755 1710
rect 5770 1410 5805 1710
rect 5975 1260 6010 1560
rect 6025 1260 6060 1560
rect 6325 1410 6360 1710
rect 6375 1410 6410 1710
rect 6990 1705 7025 1715
rect 6990 1675 6995 1705
rect 7015 1675 7025 1705
rect 6990 1640 7025 1675
rect 6990 1610 6995 1640
rect 7015 1610 7025 1640
rect 5715 930 5750 940
rect 5715 900 5720 930
rect 5740 900 5750 930
rect 5715 865 5750 900
rect 5715 835 5720 865
rect 5740 835 5750 865
rect 5715 805 5750 835
rect 5715 775 5720 805
rect 5740 775 5750 805
rect 5715 740 5750 775
rect 5715 710 5720 740
rect 5740 710 5750 740
rect 5715 680 5750 710
rect 5715 650 5720 680
rect 5740 650 5750 680
rect 5715 640 5750 650
rect 5765 930 5800 940
rect 5765 900 5775 930
rect 5795 900 5800 930
rect 5765 870 5800 900
rect 5765 840 5775 870
rect 5795 840 5800 870
rect 5765 805 5800 840
rect 5765 775 5775 805
rect 5795 775 5800 805
rect 5765 745 5800 775
rect 5765 715 5775 745
rect 5795 715 5800 745
rect 5765 680 5800 715
rect 5765 650 5775 680
rect 5795 650 5800 680
rect 5765 640 5800 650
rect 5970 780 6005 790
rect 5970 750 5975 780
rect 5995 750 6005 780
rect 5970 715 6005 750
rect 5970 685 5975 715
rect 5995 685 6005 715
rect 5970 655 6005 685
rect 5970 625 5975 655
rect 5995 625 6005 655
rect 5970 590 6005 625
rect 5970 560 5975 590
rect 5995 560 6005 590
rect 5970 530 6005 560
rect 5970 500 5975 530
rect 5995 500 6005 530
rect 5970 490 6005 500
rect 6020 780 6055 790
rect 6020 750 6030 780
rect 6050 750 6055 780
rect 6020 720 6055 750
rect 6020 690 6030 720
rect 6050 690 6055 720
rect 6020 655 6055 690
rect 6020 625 6030 655
rect 6050 625 6055 655
rect 6020 595 6055 625
rect 6020 565 6030 595
rect 6050 565 6055 595
rect 6020 530 6055 565
rect 6020 500 6030 530
rect 6050 500 6055 530
rect 6020 490 6055 500
rect 6580 1260 6615 1560
rect 6630 1260 6665 1560
rect 6990 1580 7025 1610
rect 6990 1550 6995 1580
rect 7015 1550 7025 1580
rect 6990 1515 7025 1550
rect 6990 1485 6995 1515
rect 7015 1485 7025 1515
rect 6990 1455 7025 1485
rect 6990 1425 6995 1455
rect 7015 1425 7025 1455
rect 6990 1415 7025 1425
rect 7040 1705 7075 1715
rect 7040 1675 7050 1705
rect 7070 1675 7075 1705
rect 7040 1645 7075 1675
rect 7040 1615 7050 1645
rect 7070 1615 7075 1645
rect 7585 1705 7620 1715
rect 7585 1675 7590 1705
rect 7610 1675 7620 1705
rect 7585 1640 7620 1675
rect 7040 1580 7075 1615
rect 7585 1610 7590 1640
rect 7610 1610 7620 1640
rect 7040 1550 7050 1580
rect 7070 1550 7075 1580
rect 7040 1520 7075 1550
rect 7040 1490 7050 1520
rect 7070 1490 7075 1520
rect 7040 1455 7075 1490
rect 7040 1425 7050 1455
rect 7070 1425 7075 1455
rect 7040 1415 7075 1425
rect 7245 1555 7280 1565
rect 7245 1525 7250 1555
rect 7270 1525 7280 1555
rect 7245 1490 7280 1525
rect 7245 1460 7250 1490
rect 7270 1460 7280 1490
rect 7245 1430 7280 1460
rect 6320 930 6355 940
rect 6320 900 6325 930
rect 6345 900 6355 930
rect 6320 865 6355 900
rect 6320 835 6325 865
rect 6345 835 6355 865
rect 6320 805 6355 835
rect 6320 775 6325 805
rect 6345 775 6355 805
rect 6320 740 6355 775
rect 6320 710 6325 740
rect 6345 710 6355 740
rect 6320 680 6355 710
rect 6320 650 6325 680
rect 6345 650 6355 680
rect 6320 640 6355 650
rect 6370 930 6405 940
rect 6370 900 6380 930
rect 6400 900 6405 930
rect 6370 870 6405 900
rect 6370 840 6380 870
rect 6400 840 6405 870
rect 6370 805 6405 840
rect 6370 775 6380 805
rect 6400 775 6405 805
rect 7245 1400 7250 1430
rect 7270 1400 7280 1430
rect 7245 1365 7280 1400
rect 7245 1335 7250 1365
rect 7270 1335 7280 1365
rect 7245 1305 7280 1335
rect 7245 1275 7250 1305
rect 7270 1275 7280 1305
rect 7245 1265 7280 1275
rect 7295 1555 7330 1565
rect 7295 1525 7305 1555
rect 7325 1525 7330 1555
rect 7295 1495 7330 1525
rect 7295 1465 7305 1495
rect 7325 1465 7330 1495
rect 7295 1430 7330 1465
rect 7295 1400 7305 1430
rect 7325 1400 7330 1430
rect 7295 1370 7330 1400
rect 7295 1340 7305 1370
rect 7325 1340 7330 1370
rect 7295 1305 7330 1340
rect 7295 1275 7305 1305
rect 7325 1275 7330 1305
rect 7295 1265 7330 1275
rect 7585 1580 7620 1610
rect 7585 1550 7590 1580
rect 7610 1550 7620 1580
rect 7585 1515 7620 1550
rect 7585 1485 7590 1515
rect 7610 1485 7620 1515
rect 7585 1455 7620 1485
rect 7585 1425 7590 1455
rect 7610 1425 7620 1455
rect 7585 1415 7620 1425
rect 7635 1705 7670 1715
rect 7635 1675 7645 1705
rect 7665 1675 7670 1705
rect 7635 1645 7670 1675
rect 7635 1615 7645 1645
rect 7665 1615 7670 1645
rect 7635 1580 7670 1615
rect 7635 1550 7645 1580
rect 7665 1550 7670 1580
rect 7635 1520 7670 1550
rect 7635 1490 7645 1520
rect 7665 1490 7670 1520
rect 7635 1455 7670 1490
rect 7635 1425 7645 1455
rect 7665 1425 7670 1455
rect 7635 1415 7670 1425
rect 7840 1555 7875 1565
rect 7840 1525 7845 1555
rect 7865 1525 7875 1555
rect 7840 1490 7875 1525
rect 7840 1460 7845 1490
rect 7865 1460 7875 1490
rect 7840 1430 7875 1460
rect 7840 1400 7845 1430
rect 7865 1400 7875 1430
rect 7840 1365 7875 1400
rect 7840 1335 7845 1365
rect 7865 1335 7875 1365
rect 7840 1305 7875 1335
rect 7840 1275 7845 1305
rect 7865 1275 7875 1305
rect 7840 1265 7875 1275
rect 7890 1555 7925 1565
rect 7890 1525 7900 1555
rect 7920 1525 7925 1555
rect 7890 1495 7925 1525
rect 7890 1465 7900 1495
rect 7920 1465 7925 1495
rect 7890 1430 7925 1465
rect 7890 1400 7900 1430
rect 7920 1400 7925 1430
rect 7890 1370 7925 1400
rect 7890 1340 7900 1370
rect 7920 1340 7925 1370
rect 7890 1305 7925 1340
rect 7890 1275 7900 1305
rect 7920 1275 7925 1305
rect 7890 1265 7925 1275
rect 6370 745 6405 775
rect 6370 715 6380 745
rect 6400 715 6405 745
rect 6370 680 6405 715
rect 6370 650 6380 680
rect 6400 650 6405 680
rect 6370 640 6405 650
rect 6575 780 6610 790
rect 6575 750 6580 780
rect 6600 750 6610 780
rect 6575 715 6610 750
rect 6575 685 6580 715
rect 6600 685 6610 715
rect 6575 655 6610 685
rect 6575 625 6580 655
rect 6600 625 6610 655
rect 6575 590 6610 625
rect 6575 560 6580 590
rect 6600 560 6610 590
rect 6575 530 6610 560
rect 6575 500 6580 530
rect 6600 500 6610 530
rect 6575 490 6610 500
rect 6625 780 6660 790
rect 6625 750 6635 780
rect 6655 750 6660 780
rect 6625 720 6660 750
rect 6625 690 6635 720
rect 6655 690 6660 720
rect 6625 655 6660 690
rect 6625 625 6635 655
rect 6655 625 6660 655
rect 6625 595 6660 625
rect 6625 565 6635 595
rect 6655 565 6660 595
rect 6625 530 6660 565
rect 6985 935 7020 945
rect 6985 905 6990 935
rect 7010 905 7020 935
rect 6985 870 7020 905
rect 6985 840 6990 870
rect 7010 840 7020 870
rect 6985 810 7020 840
rect 6985 780 6990 810
rect 7010 780 7020 810
rect 6985 745 7020 780
rect 6985 715 6990 745
rect 7010 715 7020 745
rect 6985 685 7020 715
rect 6985 655 6990 685
rect 7010 655 7020 685
rect 6985 645 7020 655
rect 7035 935 7070 945
rect 7035 905 7045 935
rect 7065 905 7070 935
rect 7035 875 7070 905
rect 7035 845 7045 875
rect 7065 845 7070 875
rect 7580 935 7615 945
rect 7580 905 7585 935
rect 7605 905 7615 935
rect 7580 870 7615 905
rect 7035 810 7070 845
rect 7580 840 7585 870
rect 7605 840 7615 870
rect 7580 810 7615 840
rect 7035 780 7045 810
rect 7065 780 7070 810
rect 7035 750 7070 780
rect 7035 720 7045 750
rect 7065 720 7070 750
rect 7035 685 7070 720
rect 7035 655 7045 685
rect 7065 655 7070 685
rect 7035 645 7070 655
rect 7240 785 7275 795
rect 7240 755 7245 785
rect 7265 755 7275 785
rect 7240 720 7275 755
rect 7240 690 7245 720
rect 7265 690 7275 720
rect 7240 660 7275 690
rect 7240 630 7245 660
rect 7265 630 7275 660
rect 7240 595 7275 630
rect 6625 500 6635 530
rect 6655 500 6660 530
rect 6625 490 6660 500
rect 7240 565 7245 595
rect 7265 565 7275 595
rect 7240 535 7275 565
rect 7240 505 7245 535
rect 7265 505 7275 535
rect 7240 495 7275 505
rect 7290 785 7325 795
rect 7290 755 7300 785
rect 7320 755 7325 785
rect 7290 725 7325 755
rect 7580 780 7585 810
rect 7605 780 7615 810
rect 7290 695 7300 725
rect 7320 695 7325 725
rect 7290 660 7325 695
rect 7290 630 7300 660
rect 7320 630 7325 660
rect 7290 600 7325 630
rect 7290 570 7300 600
rect 7320 570 7325 600
rect 7290 535 7325 570
rect 7290 505 7300 535
rect 7320 505 7325 535
rect 7290 495 7325 505
rect 7580 745 7615 780
rect 7580 715 7585 745
rect 7605 715 7615 745
rect 7580 685 7615 715
rect 7580 655 7585 685
rect 7605 655 7615 685
rect 7580 645 7615 655
rect 7630 935 7665 945
rect 7630 905 7640 935
rect 7660 905 7665 935
rect 7630 875 7665 905
rect 7630 845 7640 875
rect 7660 845 7665 875
rect 9220 940 9270 1525
rect 9370 1510 9420 1525
rect 9370 1480 9380 1510
rect 9410 1480 9420 1510
rect 9370 1460 9420 1480
rect 9370 1430 9380 1460
rect 9410 1430 9420 1460
rect 9370 1410 9420 1430
rect 9370 1380 9380 1410
rect 9410 1380 9420 1410
rect 9370 1360 9420 1380
rect 9370 1330 9380 1360
rect 9410 1330 9420 1360
rect 9370 1310 9420 1330
rect 9370 1280 9380 1310
rect 9410 1280 9420 1310
rect 9370 1260 9420 1280
rect 9370 1230 9380 1260
rect 9410 1230 9420 1260
rect 9370 1210 9420 1230
rect 9370 1180 9380 1210
rect 9410 1180 9420 1210
rect 9370 1160 9420 1180
rect 9370 1130 9380 1160
rect 9410 1130 9420 1160
rect 9370 1110 9420 1130
rect 9370 1080 9380 1110
rect 9410 1080 9420 1110
rect 9370 1060 9420 1080
rect 9370 1030 9380 1060
rect 9410 1030 9420 1060
rect 9370 1010 9420 1030
rect 9370 980 9380 1010
rect 9410 980 9420 1010
rect 9370 940 9420 980
rect 9520 1510 9570 1525
rect 9520 1480 9530 1510
rect 9560 1480 9570 1510
rect 9520 1460 9570 1480
rect 9520 1430 9530 1460
rect 9560 1430 9570 1460
rect 9520 1410 9570 1430
rect 9520 1380 9530 1410
rect 9560 1380 9570 1410
rect 9520 1360 9570 1380
rect 9520 1330 9530 1360
rect 9560 1330 9570 1360
rect 9520 1310 9570 1330
rect 9520 1280 9530 1310
rect 9560 1280 9570 1310
rect 9520 1260 9570 1280
rect 9520 1230 9530 1260
rect 9560 1230 9570 1260
rect 9520 1210 9570 1230
rect 9520 1180 9530 1210
rect 9560 1180 9570 1210
rect 9520 1160 9570 1180
rect 9520 1130 9530 1160
rect 9560 1130 9570 1160
rect 9520 1110 9570 1130
rect 9520 1080 9530 1110
rect 9560 1080 9570 1110
rect 9520 1060 9570 1080
rect 9520 1030 9530 1060
rect 9560 1030 9570 1060
rect 9520 1010 9570 1030
rect 9520 980 9530 1010
rect 9560 980 9570 1010
rect 9520 940 9570 980
rect 9670 1510 9820 1525
rect 9670 1480 9680 1510
rect 9710 1480 9780 1510
rect 9810 1480 9820 1510
rect 9670 1460 9820 1480
rect 9670 1430 9680 1460
rect 9710 1430 9780 1460
rect 9810 1430 9820 1460
rect 9670 1410 9820 1430
rect 9670 1380 9680 1410
rect 9710 1380 9780 1410
rect 9810 1380 9820 1410
rect 9670 1360 9820 1380
rect 9670 1330 9680 1360
rect 9710 1330 9780 1360
rect 9810 1330 9820 1360
rect 9670 1310 9820 1330
rect 9670 1280 9680 1310
rect 9710 1280 9780 1310
rect 9810 1280 9820 1310
rect 9670 1260 9820 1280
rect 9670 1230 9680 1260
rect 9710 1230 9780 1260
rect 9810 1230 9820 1260
rect 9670 1210 9820 1230
rect 9670 1180 9680 1210
rect 9710 1180 9780 1210
rect 9810 1180 9820 1210
rect 9670 1160 9820 1180
rect 9670 1130 9680 1160
rect 9710 1130 9780 1160
rect 9810 1130 9820 1160
rect 9670 1110 9820 1130
rect 9670 1080 9680 1110
rect 9710 1080 9780 1110
rect 9810 1080 9820 1110
rect 9670 1060 9820 1080
rect 9670 1030 9680 1060
rect 9710 1030 9780 1060
rect 9810 1030 9820 1060
rect 9670 1010 9820 1030
rect 9670 980 9680 1010
rect 9710 980 9780 1010
rect 9810 980 9820 1010
rect 9670 940 9820 980
rect 9920 1510 9970 1525
rect 9920 1480 9930 1510
rect 9960 1480 9970 1510
rect 9920 1460 9970 1480
rect 9920 1430 9930 1460
rect 9960 1430 9970 1460
rect 9920 1410 9970 1430
rect 9920 1380 9930 1410
rect 9960 1380 9970 1410
rect 9920 1360 9970 1380
rect 9920 1330 9930 1360
rect 9960 1330 9970 1360
rect 9920 1310 9970 1330
rect 9920 1280 9930 1310
rect 9960 1280 9970 1310
rect 9920 1260 9970 1280
rect 9920 1230 9930 1260
rect 9960 1230 9970 1260
rect 9920 1210 9970 1230
rect 9920 1180 9930 1210
rect 9960 1180 9970 1210
rect 9920 1160 9970 1180
rect 9920 1130 9930 1160
rect 9960 1130 9970 1160
rect 9920 1110 9970 1130
rect 9920 1080 9930 1110
rect 9960 1080 9970 1110
rect 9920 1060 9970 1080
rect 9920 1030 9930 1060
rect 9960 1030 9970 1060
rect 9920 1010 9970 1030
rect 9920 980 9930 1010
rect 9960 980 9970 1010
rect 9920 940 9970 980
rect 10070 1510 10120 1525
rect 10070 1480 10080 1510
rect 10110 1480 10120 1510
rect 10070 1460 10120 1480
rect 10070 1430 10080 1460
rect 10110 1430 10120 1460
rect 10070 1410 10120 1430
rect 10070 1380 10080 1410
rect 10110 1380 10120 1410
rect 10070 1360 10120 1380
rect 10070 1330 10080 1360
rect 10110 1330 10120 1360
rect 10070 1310 10120 1330
rect 10070 1280 10080 1310
rect 10110 1280 10120 1310
rect 10070 1260 10120 1280
rect 10070 1230 10080 1260
rect 10110 1230 10120 1260
rect 10070 1210 10120 1230
rect 10070 1180 10080 1210
rect 10110 1180 10120 1210
rect 10070 1160 10120 1180
rect 10070 1130 10080 1160
rect 10110 1130 10120 1160
rect 10070 1110 10120 1130
rect 10070 1080 10080 1110
rect 10110 1080 10120 1110
rect 10070 1060 10120 1080
rect 10070 1030 10080 1060
rect 10110 1030 10120 1060
rect 10070 1010 10120 1030
rect 10070 980 10080 1010
rect 10110 980 10120 1010
rect 10070 940 10120 980
rect 10220 1510 10270 1525
rect 10220 1480 10230 1510
rect 10260 1480 10270 1510
rect 10220 1460 10270 1480
rect 10220 1430 10230 1460
rect 10260 1430 10270 1460
rect 10220 1410 10270 1430
rect 10220 1380 10230 1410
rect 10260 1380 10270 1410
rect 10220 1360 10270 1380
rect 10220 1330 10230 1360
rect 10260 1330 10270 1360
rect 10220 1310 10270 1330
rect 10220 1280 10230 1310
rect 10260 1280 10270 1310
rect 10220 1260 10270 1280
rect 10220 1230 10230 1260
rect 10260 1230 10270 1260
rect 10220 1210 10270 1230
rect 10220 1180 10230 1210
rect 10260 1180 10270 1210
rect 10220 1160 10270 1180
rect 10220 1130 10230 1160
rect 10260 1130 10270 1160
rect 10220 1110 10270 1130
rect 10220 1080 10230 1110
rect 10260 1080 10270 1110
rect 10220 1060 10270 1080
rect 10220 1030 10230 1060
rect 10260 1030 10270 1060
rect 10220 1010 10270 1030
rect 10220 980 10230 1010
rect 10260 980 10270 1010
rect 10220 940 10270 980
rect 10370 1510 10420 1525
rect 10370 1480 10380 1510
rect 10410 1480 10420 1510
rect 10370 1460 10420 1480
rect 10370 1430 10380 1460
rect 10410 1430 10420 1460
rect 10370 1410 10420 1430
rect 10370 1380 10380 1410
rect 10410 1380 10420 1410
rect 10370 1360 10420 1380
rect 10370 1330 10380 1360
rect 10410 1330 10420 1360
rect 10370 1310 10420 1330
rect 10370 1280 10380 1310
rect 10410 1280 10420 1310
rect 10370 1260 10420 1280
rect 10370 1230 10380 1260
rect 10410 1230 10420 1260
rect 10370 1210 10420 1230
rect 10370 1180 10380 1210
rect 10410 1180 10420 1210
rect 10370 1160 10420 1180
rect 10370 1130 10380 1160
rect 10410 1130 10420 1160
rect 10370 1110 10420 1130
rect 10370 1080 10380 1110
rect 10410 1080 10420 1110
rect 10370 1060 10420 1080
rect 10370 1030 10380 1060
rect 10410 1030 10420 1060
rect 10370 1010 10420 1030
rect 10370 980 10380 1010
rect 10410 980 10420 1010
rect 10370 940 10420 980
rect 10520 1510 10570 1525
rect 10520 1480 10530 1510
rect 10560 1480 10570 1510
rect 10520 1460 10570 1480
rect 10520 1430 10530 1460
rect 10560 1430 10570 1460
rect 10520 1410 10570 1430
rect 10520 1380 10530 1410
rect 10560 1380 10570 1410
rect 10520 1360 10570 1380
rect 10520 1330 10530 1360
rect 10560 1330 10570 1360
rect 10520 1310 10570 1330
rect 10520 1280 10530 1310
rect 10560 1280 10570 1310
rect 10520 1260 10570 1280
rect 10520 1230 10530 1260
rect 10560 1230 10570 1260
rect 10520 1210 10570 1230
rect 10520 1180 10530 1210
rect 10560 1180 10570 1210
rect 10520 1160 10570 1180
rect 10520 1130 10530 1160
rect 10560 1130 10570 1160
rect 10520 1110 10570 1130
rect 10520 1080 10530 1110
rect 10560 1080 10570 1110
rect 10520 1060 10570 1080
rect 10520 1030 10530 1060
rect 10560 1030 10570 1060
rect 10520 1010 10570 1030
rect 10520 980 10530 1010
rect 10560 980 10570 1010
rect 10520 940 10570 980
rect 10670 1510 10720 1525
rect 10670 1480 10680 1510
rect 10710 1480 10720 1510
rect 10670 1460 10720 1480
rect 10670 1430 10680 1460
rect 10710 1430 10720 1460
rect 10670 1410 10720 1430
rect 10670 1380 10680 1410
rect 10710 1380 10720 1410
rect 10670 1360 10720 1380
rect 10670 1330 10680 1360
rect 10710 1330 10720 1360
rect 10670 1310 10720 1330
rect 10670 1280 10680 1310
rect 10710 1280 10720 1310
rect 10670 1260 10720 1280
rect 10670 1230 10680 1260
rect 10710 1230 10720 1260
rect 10670 1210 10720 1230
rect 10670 1180 10680 1210
rect 10710 1180 10720 1210
rect 10670 1160 10720 1180
rect 10670 1130 10680 1160
rect 10710 1130 10720 1160
rect 10670 1110 10720 1130
rect 10670 1080 10680 1110
rect 10710 1080 10720 1110
rect 10670 1060 10720 1080
rect 10670 1030 10680 1060
rect 10710 1030 10720 1060
rect 10670 1010 10720 1030
rect 10670 980 10680 1010
rect 10710 980 10720 1010
rect 10670 940 10720 980
rect 10820 940 10870 1525
rect 7630 810 7665 845
rect 7630 780 7640 810
rect 7660 780 7665 810
rect 7630 750 7665 780
rect 7630 720 7640 750
rect 7660 720 7665 750
rect 7630 685 7665 720
rect 7630 655 7640 685
rect 7660 655 7665 685
rect 7630 645 7665 655
rect 7835 785 7870 795
rect 7835 755 7840 785
rect 7860 755 7870 785
rect 7835 720 7870 755
rect 7835 690 7840 720
rect 7860 690 7870 720
rect 7835 660 7870 690
rect 7835 630 7840 660
rect 7860 630 7870 660
rect 7835 595 7870 630
rect 5225 -320 5260 -20
rect 5275 -320 5310 -20
rect 5715 -170 5750 130
rect 5765 -170 5800 130
rect 7835 565 7840 595
rect 7860 565 7870 595
rect 7835 535 7870 565
rect 7835 505 7840 535
rect 7860 505 7870 535
rect 7835 495 7870 505
rect 7885 785 7920 795
rect 7885 755 7895 785
rect 7915 755 7920 785
rect 7885 725 7920 755
rect 7885 695 7895 725
rect 7915 695 7920 725
rect 7885 660 7920 695
rect 7885 630 7895 660
rect 7915 630 7920 660
rect 7885 600 7920 630
rect 7885 570 7895 600
rect 7915 570 7920 600
rect 7885 535 7920 570
rect 7885 505 7895 535
rect 7915 505 7920 535
rect 7885 495 7920 505
rect 9220 380 9270 673
rect 9370 660 9420 673
rect 9370 630 9380 660
rect 9410 630 9420 660
rect 9370 610 9420 630
rect 9370 580 9380 610
rect 9410 580 9420 610
rect 9370 560 9420 580
rect 9370 530 9380 560
rect 9410 530 9420 560
rect 9370 510 9420 530
rect 9370 480 9380 510
rect 9410 480 9420 510
rect 9370 460 9420 480
rect 9370 400 9380 460
rect 9410 400 9420 460
rect 9370 380 9420 400
rect 9520 660 9570 673
rect 9520 630 9530 660
rect 9560 630 9570 660
rect 9520 610 9570 630
rect 9520 580 9530 610
rect 9560 580 9570 610
rect 9520 560 9570 580
rect 9520 530 9530 560
rect 9560 530 9570 560
rect 9520 510 9570 530
rect 9520 480 9530 510
rect 9560 480 9570 510
rect 9520 460 9570 480
rect 9520 400 9530 460
rect 9560 400 9570 460
rect 9520 380 9570 400
rect 9670 660 9720 673
rect 9670 630 9680 660
rect 9710 630 9720 660
rect 9670 610 9720 630
rect 9670 580 9680 610
rect 9710 580 9720 610
rect 9670 560 9720 580
rect 9670 530 9680 560
rect 9710 530 9720 560
rect 9670 510 9720 530
rect 9670 480 9680 510
rect 9710 480 9720 510
rect 9670 460 9720 480
rect 9670 400 9680 460
rect 9710 400 9720 460
rect 9670 380 9720 400
rect 9820 380 9870 673
rect 5970 -320 6005 -20
rect 6020 -320 6055 -20
rect 6320 -170 6355 130
rect 6370 -170 6405 130
rect 6575 -320 6610 -20
rect 6625 -320 6660 -20
rect 6985 -165 7020 135
rect 7035 -165 7070 135
rect 7580 125 7615 135
rect 7580 95 7585 125
rect 7605 95 7615 125
rect 7580 60 7615 95
rect 7580 30 7585 60
rect 7605 30 7615 60
rect 7580 0 7615 30
rect 7240 -315 7275 -15
rect 7290 -315 7325 -15
rect 7580 -30 7585 0
rect 7605 -30 7615 0
rect 7580 -65 7615 -30
rect 7580 -95 7585 -65
rect 7605 -95 7615 -65
rect 7580 -125 7615 -95
rect 7580 -155 7585 -125
rect 7605 -155 7615 -125
rect 7580 -165 7615 -155
rect 7630 125 7665 135
rect 7630 95 7640 125
rect 7660 95 7665 125
rect 7630 65 7665 95
rect 7630 35 7640 65
rect 7660 35 7665 65
rect 7630 0 7665 35
rect 7630 -30 7640 0
rect 7660 -30 7665 0
rect 7630 -60 7665 -30
rect 7630 -90 7640 -60
rect 7660 -90 7665 -60
rect 7630 -125 7665 -90
rect 7630 -155 7640 -125
rect 7660 -155 7665 -125
rect 7630 -165 7665 -155
rect 7835 -25 7870 -15
rect 7835 -55 7840 -25
rect 7860 -55 7870 -25
rect 7835 -90 7870 -55
rect 7835 -120 7840 -90
rect 7860 -120 7870 -90
rect 7835 -150 7870 -120
rect 7835 -180 7840 -150
rect 7860 -180 7870 -150
rect 7835 -215 7870 -180
rect 7835 -245 7840 -215
rect 7860 -245 7870 -215
rect 7835 -275 7870 -245
rect 7835 -305 7840 -275
rect 7860 -305 7870 -275
rect 7835 -315 7870 -305
rect 7885 -25 7920 -15
rect 7885 -55 7895 -25
rect 7915 -55 7920 -25
rect 7885 -85 7920 -55
rect 7885 -115 7895 -85
rect 7915 -115 7920 -85
rect 7885 -150 7920 -115
rect 7885 -180 7895 -150
rect 7915 -180 7920 -150
rect 7885 -210 7920 -180
rect 7885 -240 7895 -210
rect 7915 -240 7920 -210
rect 7885 -275 7920 -240
rect 7885 -305 7895 -275
rect 7915 -305 7920 -275
rect 7885 -315 7920 -305
rect 10590 41 10620 626
rect 10720 590 10770 626
rect 10720 560 10730 590
rect 10760 560 10770 590
rect 10720 540 10770 560
rect 10720 510 10730 540
rect 10760 510 10770 540
rect 10720 490 10770 510
rect 10720 460 10730 490
rect 10760 460 10770 490
rect 10720 440 10770 460
rect 10720 410 10730 440
rect 10760 410 10770 440
rect 10720 390 10770 410
rect 10720 360 10730 390
rect 10760 360 10770 390
rect 10720 340 10770 360
rect 10720 310 10730 340
rect 10760 310 10770 340
rect 10720 290 10770 310
rect 10720 260 10730 290
rect 10760 260 10770 290
rect 10720 240 10770 260
rect 10720 210 10730 240
rect 10760 210 10770 240
rect 10720 190 10770 210
rect 10720 160 10730 190
rect 10760 160 10770 190
rect 10720 140 10770 160
rect 10720 110 10730 140
rect 10760 110 10770 140
rect 10720 90 10770 110
rect 10720 60 10730 90
rect 10760 60 10770 90
rect 10720 41 10770 60
rect 10870 590 10920 626
rect 10870 560 10880 590
rect 10910 560 10920 590
rect 10870 540 10920 560
rect 10870 510 10880 540
rect 10910 510 10920 540
rect 10870 490 10920 510
rect 10870 460 10880 490
rect 10910 460 10920 490
rect 10870 440 10920 460
rect 10870 410 10880 440
rect 10910 410 10920 440
rect 10870 390 10920 410
rect 10870 360 10880 390
rect 10910 360 10920 390
rect 10870 340 10920 360
rect 10870 310 10880 340
rect 10910 310 10920 340
rect 10870 290 10920 310
rect 10870 260 10880 290
rect 10910 260 10920 290
rect 10870 240 10920 260
rect 10870 210 10880 240
rect 10910 210 10920 240
rect 10870 190 10920 210
rect 10870 160 10880 190
rect 10910 160 10920 190
rect 10870 140 10920 160
rect 10870 110 10880 140
rect 10910 110 10920 140
rect 10870 90 10920 110
rect 10870 60 10880 90
rect 10910 60 10920 90
rect 10870 41 10920 60
rect 11020 41 11050 626
<< ndiffc >>
rect 5230 910 5250 940
rect 5230 860 5250 890
rect 5285 910 5305 940
rect 5285 860 5305 890
rect 4975 525 4995 555
rect 4975 475 4995 505
rect 5030 525 5050 555
rect 5030 475 5050 505
rect 5975 910 5995 940
rect 5975 860 5995 890
rect 6030 910 6050 940
rect 6030 860 6050 890
rect 5720 525 5740 555
rect 5720 475 5740 505
rect 5775 525 5795 555
rect 5775 475 5795 505
rect 7250 1685 7270 1715
rect 7250 1635 7270 1665
rect 7305 1685 7325 1715
rect 7305 1635 7325 1665
rect 6580 910 6600 940
rect 6580 860 6600 890
rect 6635 910 6655 940
rect 6635 860 6655 890
rect 6995 1300 7015 1330
rect 6995 1250 7015 1280
rect 7050 1300 7070 1330
rect 7050 1250 7070 1280
rect 7845 1685 7865 1715
rect 7845 1635 7865 1665
rect 7900 1685 7920 1715
rect 7900 1635 7920 1665
rect 7590 1300 7610 1330
rect 7590 1250 7610 1280
rect 7645 1300 7665 1330
rect 7645 1250 7665 1280
rect 6325 525 6345 555
rect 6325 475 6345 505
rect 6380 525 6400 555
rect 6380 475 6400 505
rect 7245 915 7265 945
rect 7245 865 7265 895
rect 7300 915 7320 945
rect 7300 865 7320 895
rect 6990 530 7010 560
rect 6990 480 7010 510
rect 7045 530 7065 560
rect 7045 480 7065 510
rect 7840 915 7860 945
rect 7840 865 7860 895
rect 7895 915 7915 945
rect 7895 865 7915 895
rect 7585 530 7605 560
rect 7585 480 7605 510
rect 7640 530 7660 560
rect 7640 480 7660 510
rect 7840 105 7860 135
rect 7840 55 7860 85
rect 7895 105 7915 135
rect 7895 55 7915 85
rect 7585 -280 7605 -250
rect 7585 -330 7605 -300
rect 7640 -280 7660 -250
rect 7640 -330 7660 -300
rect 9380 -50 9410 0
rect 9530 -50 9560 0
rect 9680 -50 9710 0
rect 10150 600 10180 630
rect 10150 550 10180 580
rect 10150 500 10180 530
rect 10150 450 10180 480
rect 10150 400 10180 430
rect 10150 350 10180 380
rect 10150 300 10180 330
rect 10150 250 10180 280
rect 10150 200 10180 230
rect 10150 150 10180 180
rect 10150 100 10180 130
rect 10150 50 10180 80
rect 10150 0 10180 30
rect 10150 -50 10180 -20
rect 10150 -100 10180 -70
rect 10150 -150 10180 -120
rect 10150 -200 10180 -170
rect 10300 600 10330 630
rect 10300 550 10330 580
rect 10300 500 10330 530
rect 10300 450 10330 480
rect 10300 400 10330 430
rect 10300 350 10330 380
rect 10300 300 10330 330
rect 10300 250 10330 280
rect 10300 200 10330 230
rect 10300 150 10330 180
rect 10300 100 10330 130
rect 10300 50 10330 80
rect 10300 0 10330 30
rect 10300 -50 10330 -20
rect 10300 -100 10330 -70
rect 10300 -150 10330 -120
rect 10300 -200 10330 -170
<< pdiffc >>
rect 4975 900 4995 930
rect 4975 835 4995 865
rect 4975 775 4995 805
rect 4975 710 4995 740
rect 4975 650 4995 680
rect 5030 900 5050 930
rect 5030 840 5050 870
rect 5030 775 5050 805
rect 5030 715 5050 745
rect 5030 650 5050 680
rect 5230 750 5250 780
rect 5230 685 5250 715
rect 5230 625 5250 655
rect 5230 560 5250 590
rect 5230 500 5250 530
rect 5285 750 5305 780
rect 5285 690 5305 720
rect 5285 625 5305 655
rect 5285 565 5305 595
rect 5285 500 5305 530
rect 6995 1675 7015 1705
rect 6995 1610 7015 1640
rect 5720 900 5740 930
rect 5720 835 5740 865
rect 5720 775 5740 805
rect 5720 710 5740 740
rect 5720 650 5740 680
rect 5775 900 5795 930
rect 5775 840 5795 870
rect 5775 775 5795 805
rect 5775 715 5795 745
rect 5775 650 5795 680
rect 5975 750 5995 780
rect 5975 685 5995 715
rect 5975 625 5995 655
rect 5975 560 5995 590
rect 5975 500 5995 530
rect 6030 750 6050 780
rect 6030 690 6050 720
rect 6030 625 6050 655
rect 6030 565 6050 595
rect 6030 500 6050 530
rect 6995 1550 7015 1580
rect 6995 1485 7015 1515
rect 6995 1425 7015 1455
rect 7050 1675 7070 1705
rect 7050 1615 7070 1645
rect 7590 1675 7610 1705
rect 7590 1610 7610 1640
rect 7050 1550 7070 1580
rect 7050 1490 7070 1520
rect 7050 1425 7070 1455
rect 7250 1525 7270 1555
rect 7250 1460 7270 1490
rect 6325 900 6345 930
rect 6325 835 6345 865
rect 6325 775 6345 805
rect 6325 710 6345 740
rect 6325 650 6345 680
rect 6380 900 6400 930
rect 6380 840 6400 870
rect 6380 775 6400 805
rect 7250 1400 7270 1430
rect 7250 1335 7270 1365
rect 7250 1275 7270 1305
rect 7305 1525 7325 1555
rect 7305 1465 7325 1495
rect 7305 1400 7325 1430
rect 7305 1340 7325 1370
rect 7305 1275 7325 1305
rect 7590 1550 7610 1580
rect 7590 1485 7610 1515
rect 7590 1425 7610 1455
rect 7645 1675 7665 1705
rect 7645 1615 7665 1645
rect 7645 1550 7665 1580
rect 7645 1490 7665 1520
rect 7645 1425 7665 1455
rect 7845 1525 7865 1555
rect 7845 1460 7865 1490
rect 7845 1400 7865 1430
rect 7845 1335 7865 1365
rect 7845 1275 7865 1305
rect 7900 1525 7920 1555
rect 7900 1465 7920 1495
rect 7900 1400 7920 1430
rect 7900 1340 7920 1370
rect 7900 1275 7920 1305
rect 6380 715 6400 745
rect 6380 650 6400 680
rect 6580 750 6600 780
rect 6580 685 6600 715
rect 6580 625 6600 655
rect 6580 560 6600 590
rect 6580 500 6600 530
rect 6635 750 6655 780
rect 6635 690 6655 720
rect 6635 625 6655 655
rect 6635 565 6655 595
rect 6990 905 7010 935
rect 6990 840 7010 870
rect 6990 780 7010 810
rect 6990 715 7010 745
rect 6990 655 7010 685
rect 7045 905 7065 935
rect 7045 845 7065 875
rect 7585 905 7605 935
rect 7585 840 7605 870
rect 7045 780 7065 810
rect 7045 720 7065 750
rect 7045 655 7065 685
rect 7245 755 7265 785
rect 7245 690 7265 720
rect 7245 630 7265 660
rect 6635 500 6655 530
rect 7245 565 7265 595
rect 7245 505 7265 535
rect 7300 755 7320 785
rect 7585 780 7605 810
rect 7300 695 7320 725
rect 7300 630 7320 660
rect 7300 570 7320 600
rect 7300 505 7320 535
rect 7585 715 7605 745
rect 7585 655 7605 685
rect 7640 905 7660 935
rect 7640 845 7660 875
rect 9380 1480 9410 1510
rect 9380 1430 9410 1460
rect 9380 1380 9410 1410
rect 9380 1330 9410 1360
rect 9380 1280 9410 1310
rect 9380 1230 9410 1260
rect 9380 1180 9410 1210
rect 9380 1130 9410 1160
rect 9380 1080 9410 1110
rect 9380 1030 9410 1060
rect 9380 980 9410 1010
rect 9530 1480 9560 1510
rect 9530 1430 9560 1460
rect 9530 1380 9560 1410
rect 9530 1330 9560 1360
rect 9530 1280 9560 1310
rect 9530 1230 9560 1260
rect 9530 1180 9560 1210
rect 9530 1130 9560 1160
rect 9530 1080 9560 1110
rect 9530 1030 9560 1060
rect 9530 980 9560 1010
rect 9680 1480 9710 1510
rect 9780 1480 9810 1510
rect 9680 1430 9710 1460
rect 9780 1430 9810 1460
rect 9680 1380 9710 1410
rect 9780 1380 9810 1410
rect 9680 1330 9710 1360
rect 9780 1330 9810 1360
rect 9680 1280 9710 1310
rect 9780 1280 9810 1310
rect 9680 1230 9710 1260
rect 9780 1230 9810 1260
rect 9680 1180 9710 1210
rect 9780 1180 9810 1210
rect 9680 1130 9710 1160
rect 9780 1130 9810 1160
rect 9680 1080 9710 1110
rect 9780 1080 9810 1110
rect 9680 1030 9710 1060
rect 9780 1030 9810 1060
rect 9680 980 9710 1010
rect 9780 980 9810 1010
rect 9930 1480 9960 1510
rect 9930 1430 9960 1460
rect 9930 1380 9960 1410
rect 9930 1330 9960 1360
rect 9930 1280 9960 1310
rect 9930 1230 9960 1260
rect 9930 1180 9960 1210
rect 9930 1130 9960 1160
rect 9930 1080 9960 1110
rect 9930 1030 9960 1060
rect 9930 980 9960 1010
rect 10080 1480 10110 1510
rect 10080 1430 10110 1460
rect 10080 1380 10110 1410
rect 10080 1330 10110 1360
rect 10080 1280 10110 1310
rect 10080 1230 10110 1260
rect 10080 1180 10110 1210
rect 10080 1130 10110 1160
rect 10080 1080 10110 1110
rect 10080 1030 10110 1060
rect 10080 980 10110 1010
rect 10230 1480 10260 1510
rect 10230 1430 10260 1460
rect 10230 1380 10260 1410
rect 10230 1330 10260 1360
rect 10230 1280 10260 1310
rect 10230 1230 10260 1260
rect 10230 1180 10260 1210
rect 10230 1130 10260 1160
rect 10230 1080 10260 1110
rect 10230 1030 10260 1060
rect 10230 980 10260 1010
rect 10380 1480 10410 1510
rect 10380 1430 10410 1460
rect 10380 1380 10410 1410
rect 10380 1330 10410 1360
rect 10380 1280 10410 1310
rect 10380 1230 10410 1260
rect 10380 1180 10410 1210
rect 10380 1130 10410 1160
rect 10380 1080 10410 1110
rect 10380 1030 10410 1060
rect 10380 980 10410 1010
rect 10530 1480 10560 1510
rect 10530 1430 10560 1460
rect 10530 1380 10560 1410
rect 10530 1330 10560 1360
rect 10530 1280 10560 1310
rect 10530 1230 10560 1260
rect 10530 1180 10560 1210
rect 10530 1130 10560 1160
rect 10530 1080 10560 1110
rect 10530 1030 10560 1060
rect 10530 980 10560 1010
rect 10680 1480 10710 1510
rect 10680 1430 10710 1460
rect 10680 1380 10710 1410
rect 10680 1330 10710 1360
rect 10680 1280 10710 1310
rect 10680 1230 10710 1260
rect 10680 1180 10710 1210
rect 10680 1130 10710 1160
rect 10680 1080 10710 1110
rect 10680 1030 10710 1060
rect 10680 980 10710 1010
rect 7640 780 7660 810
rect 7640 720 7660 750
rect 7640 655 7660 685
rect 7840 755 7860 785
rect 7840 690 7860 720
rect 7840 630 7860 660
rect 7840 565 7860 595
rect 7840 505 7860 535
rect 7895 755 7915 785
rect 7895 695 7915 725
rect 7895 630 7915 660
rect 7895 570 7915 600
rect 7895 505 7915 535
rect 9380 630 9410 660
rect 9380 580 9410 610
rect 9380 530 9410 560
rect 9380 480 9410 510
rect 9380 400 9410 460
rect 9530 630 9560 660
rect 9530 580 9560 610
rect 9530 530 9560 560
rect 9530 480 9560 510
rect 9530 400 9560 460
rect 9680 630 9710 660
rect 9680 580 9710 610
rect 9680 530 9710 560
rect 9680 480 9710 510
rect 9680 400 9710 460
rect 7585 95 7605 125
rect 7585 30 7605 60
rect 7585 -30 7605 0
rect 7585 -95 7605 -65
rect 7585 -155 7605 -125
rect 7640 95 7660 125
rect 7640 35 7660 65
rect 7640 -30 7660 0
rect 7640 -90 7660 -60
rect 7640 -155 7660 -125
rect 7840 -55 7860 -25
rect 7840 -120 7860 -90
rect 7840 -180 7860 -150
rect 7840 -245 7860 -215
rect 7840 -305 7860 -275
rect 7895 -55 7915 -25
rect 7895 -115 7915 -85
rect 7895 -180 7915 -150
rect 7895 -240 7915 -210
rect 7895 -305 7915 -275
rect 10730 560 10760 590
rect 10730 510 10760 540
rect 10730 460 10760 490
rect 10730 410 10760 440
rect 10730 360 10760 390
rect 10730 310 10760 340
rect 10730 260 10760 290
rect 10730 210 10760 240
rect 10730 160 10760 190
rect 10730 110 10760 140
rect 10730 60 10760 90
rect 10880 560 10910 590
rect 10880 510 10910 540
rect 10880 460 10910 490
rect 10880 410 10910 440
rect 10880 360 10910 390
rect 10880 310 10910 340
rect 10880 260 10910 290
rect 10880 210 10910 240
rect 10880 160 10910 190
rect 10880 110 10910 140
rect 10880 60 10910 90
<< psubdiff >>
rect 10950 -200 11045 -180
rect 10950 -260 10965 -200
rect 11020 -260 11045 -200
rect 10950 -280 11045 -260
<< nsubdiff >>
rect 7030 1790 7080 1805
rect 7625 1790 7675 1805
rect 5010 1015 5060 1030
rect 5010 990 5020 1015
rect 5045 990 5060 1015
rect 5010 975 5060 990
rect 7030 1765 7040 1790
rect 7065 1765 7080 1790
rect 7030 1750 7080 1765
rect 7625 1765 7635 1790
rect 7660 1765 7675 1790
rect 7625 1750 7675 1765
rect 5755 1015 5805 1030
rect 5755 990 5765 1015
rect 5790 990 5805 1015
rect 5755 975 5805 990
rect 10580 1730 10670 1750
rect 6360 1015 6410 1030
rect 6360 990 6370 1015
rect 6395 990 6410 1015
rect 6360 975 6410 990
rect 10580 1670 10600 1730
rect 10650 1670 10670 1730
rect 10580 1650 10670 1670
rect 7025 1020 7075 1035
rect 7025 995 7035 1020
rect 7060 995 7075 1020
rect 7025 980 7075 995
rect 7620 1020 7670 1035
rect 7620 995 7630 1020
rect 7655 995 7670 1020
rect 7620 980 7670 995
rect 7620 210 7670 225
rect 7620 185 7630 210
rect 7655 185 7670 210
rect 7620 170 7670 185
<< psubdiffcont >>
rect 10965 -260 11020 -200
<< nsubdiffcont >>
rect 5020 990 5045 1015
rect 7040 1765 7065 1790
rect 7635 1765 7660 1790
rect 5765 990 5790 1015
rect 6370 990 6395 1015
rect 10600 1670 10650 1730
rect 7035 995 7060 1020
rect 7630 995 7655 1020
rect 7630 185 7655 210
<< poly >>
rect 5245 1785 5285 1825
rect 5990 1785 6030 1825
rect 6595 1785 6635 1825
rect 7260 1820 7300 1830
rect 7260 1800 7270 1820
rect 7290 1800 7300 1820
rect 7855 1820 7895 1830
rect 7260 1790 7300 1800
rect 7855 1800 7865 1820
rect 7885 1800 7895 1820
rect 7855 1790 7895 1800
rect 5010 1710 5025 1725
rect 5265 1720 5280 1785
rect 5755 1710 5770 1725
rect 6010 1720 6025 1785
rect 5265 1605 5280 1620
rect 5265 1560 5280 1575
rect 4920 1375 4960 1385
rect 5010 1375 5025 1410
rect 4920 1360 5025 1375
rect 4920 1345 4960 1360
rect 5010 1335 5025 1360
rect 5010 1220 5025 1235
rect 5265 1220 5280 1260
rect 5255 1180 5295 1220
rect 5240 1045 5280 1055
rect 5240 1025 5250 1045
rect 5270 1025 5280 1045
rect 5240 1015 5280 1025
rect 5005 940 5020 955
rect 5260 950 5275 1015
rect 5260 835 5275 850
rect 5260 790 5275 805
rect 4915 605 4955 615
rect 5005 605 5020 640
rect 4915 585 4925 605
rect 4945 590 5020 605
rect 4945 585 4955 590
rect 4915 575 4955 585
rect 5005 565 5020 590
rect 5005 450 5020 465
rect 5260 450 5275 490
rect 5250 440 5290 450
rect 5250 420 5260 440
rect 5280 420 5290 440
rect 5250 410 5290 420
rect 5240 205 5280 245
rect 5005 130 5020 145
rect 5260 140 5275 205
rect 5260 25 5275 40
rect 6360 1710 6375 1725
rect 6615 1720 6630 1785
rect 6010 1605 6025 1620
rect 6010 1560 6025 1575
rect 5665 1375 5705 1385
rect 5755 1375 5770 1410
rect 5665 1360 5770 1375
rect 5665 1345 5705 1360
rect 5755 1335 5770 1360
rect 7025 1715 7040 1730
rect 7280 1725 7295 1790
rect 6615 1605 6630 1620
rect 6615 1560 6630 1575
rect 5755 1220 5770 1235
rect 6010 1220 6025 1260
rect 6000 1180 6040 1220
rect 5985 1045 6025 1055
rect 5985 1025 5995 1045
rect 6015 1025 6025 1045
rect 5985 1015 6025 1025
rect 5750 940 5765 955
rect 6005 950 6020 1015
rect 6005 835 6020 850
rect 6005 790 6020 805
rect 5665 605 5705 615
rect 5750 605 5765 640
rect 5665 585 5675 605
rect 5695 590 5765 605
rect 5695 585 5705 590
rect 5665 575 5705 585
rect 5750 565 5765 590
rect 5750 450 5765 465
rect 6005 450 6020 490
rect 5995 440 6035 450
rect 5995 420 6005 440
rect 6025 420 6035 440
rect 5995 410 6035 420
rect 5985 205 6025 245
rect 6270 1375 6310 1385
rect 6360 1375 6375 1410
rect 6270 1360 6375 1375
rect 6270 1345 6310 1360
rect 6360 1335 6375 1360
rect 7620 1715 7635 1730
rect 7875 1725 7890 1790
rect 7280 1610 7295 1625
rect 7280 1565 7295 1580
rect 6360 1220 6375 1235
rect 6615 1220 6630 1260
rect 6605 1180 6645 1220
rect 6590 1045 6630 1055
rect 6590 1025 6600 1045
rect 6620 1025 6630 1045
rect 6590 1015 6630 1025
rect 6355 940 6370 955
rect 6610 950 6625 1015
rect 6610 835 6625 850
rect 6610 790 6625 805
rect 6935 1380 6975 1390
rect 7025 1380 7040 1415
rect 6935 1360 6945 1380
rect 6965 1365 7040 1380
rect 6965 1360 6975 1365
rect 6935 1350 6975 1360
rect 7025 1340 7040 1365
rect 7875 1610 7890 1625
rect 7875 1565 7890 1580
rect 7025 1225 7040 1240
rect 7280 1225 7295 1265
rect 7270 1215 7310 1225
rect 7270 1195 7280 1215
rect 7300 1195 7310 1215
rect 7270 1185 7310 1195
rect 7530 1380 7570 1390
rect 7620 1380 7635 1415
rect 7530 1360 7540 1380
rect 7560 1365 7635 1380
rect 7560 1360 7570 1365
rect 7530 1350 7570 1360
rect 7620 1340 7635 1365
rect 9270 1525 9370 1560
rect 9420 1525 9520 1560
rect 9570 1525 9670 1560
rect 9820 1525 9920 1560
rect 9970 1525 10070 1560
rect 10120 1525 10220 1560
rect 10270 1525 10370 1560
rect 10420 1525 10520 1560
rect 10570 1525 10670 1560
rect 10720 1525 10820 1560
rect 7620 1225 7635 1240
rect 7875 1225 7890 1265
rect 7255 1050 7295 1060
rect 7255 1030 7265 1050
rect 7285 1030 7295 1050
rect 7255 1020 7295 1030
rect 7020 945 7035 960
rect 7275 955 7290 1020
rect 7865 1215 7905 1225
rect 7865 1195 7875 1215
rect 7895 1195 7905 1215
rect 7865 1185 7905 1195
rect 7850 1050 7890 1060
rect 7850 1030 7860 1050
rect 7880 1030 7890 1050
rect 7850 1020 7890 1030
rect 6265 605 6305 615
rect 6355 605 6370 640
rect 6265 585 6275 605
rect 6295 590 6370 605
rect 6295 585 6305 590
rect 6265 575 6305 585
rect 6355 565 6370 590
rect 7615 945 7630 960
rect 7870 955 7885 1020
rect 7275 840 7290 855
rect 7275 795 7290 810
rect 6930 610 6970 620
rect 7020 610 7035 645
rect 6930 590 6940 610
rect 6960 595 7035 610
rect 6960 590 6970 595
rect 6930 580 6970 590
rect 7020 570 7035 595
rect 6355 450 6370 465
rect 6610 450 6625 490
rect 9270 920 9370 940
rect 9420 920 9520 940
rect 9570 920 9670 940
rect 9820 920 9920 940
rect 9970 920 10070 940
rect 10120 920 10220 940
rect 10270 920 10370 940
rect 10420 920 10520 940
rect 10570 920 10670 940
rect 9420 910 10670 920
rect 7870 840 7885 855
rect 7870 795 7885 810
rect 7525 610 7565 620
rect 7615 610 7630 645
rect 7525 590 7535 610
rect 7555 595 7630 610
rect 7555 590 7565 595
rect 7525 580 7565 590
rect 7615 570 7630 595
rect 7020 455 7035 470
rect 7275 455 7290 495
rect 6600 440 6640 450
rect 6600 420 6610 440
rect 6630 420 6640 440
rect 6600 410 6640 420
rect 7265 445 7305 455
rect 7265 425 7275 445
rect 7295 425 7305 445
rect 7265 415 7305 425
rect 5750 130 5765 145
rect 6005 140 6020 205
rect 5260 -20 5275 -5
rect 4915 -205 4955 -195
rect 5005 -205 5020 -170
rect 4915 -220 5020 -205
rect 4915 -235 4955 -220
rect 5005 -245 5020 -220
rect 6005 25 6020 40
rect 6590 205 6630 245
rect 7255 210 7295 250
rect 9420 870 9430 910
rect 9460 870 10670 910
rect 10720 890 10820 940
rect 7615 455 7630 470
rect 7870 455 7885 495
rect 7860 445 7900 455
rect 7860 425 7870 445
rect 7890 425 7900 445
rect 7860 415 7900 425
rect 9420 860 10670 870
rect 9270 673 9370 690
rect 9420 673 9520 690
rect 9570 673 9670 690
rect 9720 673 9820 690
rect 10040 651 10140 670
rect 10190 651 10290 670
rect 10340 651 10440 670
rect 9270 360 9370 380
rect 9030 340 9140 350
rect 9030 260 9040 340
rect 9130 330 9140 340
rect 9420 330 9520 380
rect 9130 270 9520 330
rect 9130 260 9140 270
rect 9030 250 9140 260
rect 6355 130 6370 145
rect 6610 140 6625 205
rect 6005 -20 6020 -5
rect 5660 -205 5700 -195
rect 5750 -205 5765 -170
rect 5660 -220 5765 -205
rect 5660 -235 5700 -220
rect 5750 -245 5765 -220
rect 5005 -360 5020 -345
rect 5260 -360 5275 -320
rect 7020 135 7035 150
rect 7275 145 7290 210
rect 6610 25 6625 40
rect 6610 -20 6625 -5
rect 6265 -205 6305 -195
rect 6355 -205 6370 -170
rect 6265 -220 6370 -205
rect 6265 -235 6305 -220
rect 6355 -245 6370 -220
rect 5750 -360 5765 -345
rect 6005 -360 6020 -320
rect 7275 30 7290 45
rect 7275 -15 7290 0
rect 7850 240 7890 250
rect 7850 220 7860 240
rect 7880 220 7890 240
rect 7850 210 7890 220
rect 7615 135 7630 150
rect 7870 145 7885 210
rect 9030 205 9140 220
rect 6930 -200 6970 -190
rect 7020 -200 7035 -165
rect 6930 -215 7035 -200
rect 6930 -230 6970 -215
rect 7020 -240 7035 -215
rect 6355 -360 6370 -345
rect 6610 -360 6625 -320
rect 7870 30 7885 45
rect 7870 -15 7885 0
rect 7525 -200 7565 -190
rect 7615 -200 7630 -165
rect 7525 -220 7535 -200
rect 7555 -215 7630 -200
rect 7555 -220 7565 -215
rect 7525 -230 7565 -220
rect 7615 -240 7630 -215
rect 7020 -355 7035 -340
rect 7275 -355 7290 -315
rect 9030 130 9040 205
rect 9130 200 9140 205
rect 9570 200 9670 380
rect 9720 360 9820 380
rect 9130 140 9670 200
rect 9130 130 9140 140
rect 9030 120 9140 130
rect 9420 80 9500 90
rect 9420 40 9430 80
rect 9490 40 9500 80
rect 9270 16 9370 40
rect 9420 30 9500 40
rect 9420 16 9520 30
rect 9570 16 9670 40
rect 9720 16 9820 40
rect 9270 -90 9370 -70
rect 9420 -90 9520 -70
rect 9570 -90 9670 -70
rect 9720 -90 9820 -70
rect 10620 626 10720 651
rect 10770 626 10870 651
rect 10920 626 11020 651
rect 10620 21 10720 41
rect 10770 20 10870 41
rect 10920 21 11020 41
rect 10770 10 10850 20
rect 10770 -30 10780 10
rect 10840 -30 10850 10
rect 10770 -40 10850 -30
rect 10040 -230 10140 -210
rect 10190 -230 10290 -210
rect 10340 -230 10440 -210
rect 10190 -240 10270 -230
rect 10190 -280 10210 -240
rect 10250 -280 10270 -240
rect 10190 -290 10270 -280
rect 7615 -355 7630 -340
rect 7870 -355 7885 -315
rect 5250 -400 5290 -360
rect 5995 -400 6035 -360
rect 6600 -400 6640 -360
rect 7265 -395 7305 -355
rect 7860 -365 7900 -355
rect 7860 -385 7870 -365
rect 7890 -385 7900 -365
rect 7860 -395 7900 -385
<< polycont >>
rect 7270 1800 7290 1820
rect 7865 1800 7885 1820
rect 5250 1025 5270 1045
rect 4925 585 4945 605
rect 5260 420 5280 440
rect 5995 1025 6015 1045
rect 5675 585 5695 605
rect 6005 420 6025 440
rect 6600 1025 6620 1045
rect 6945 1360 6965 1380
rect 7280 1195 7300 1215
rect 7540 1360 7560 1380
rect 7265 1030 7285 1050
rect 7875 1195 7895 1215
rect 7860 1030 7880 1050
rect 6275 585 6295 605
rect 6940 590 6960 610
rect 7535 590 7555 610
rect 6610 420 6630 440
rect 7275 425 7295 445
rect 9430 870 9460 910
rect 7870 425 7890 445
rect 9040 260 9130 340
rect 7860 220 7880 240
rect 7535 -220 7555 -200
rect 9040 130 9130 205
rect 9430 40 9490 80
rect 10780 -30 10840 10
rect 10210 -280 10250 -240
rect 7870 -385 7890 -365
<< xpolycontact >>
rect 5405 1360 5440 1600
rect 5405 0 5440 240
rect 5565 1360 5600 1600
rect 6140 1360 6175 1600
rect 5565 0 5600 240
rect 6845 1360 6880 1600
rect 7440 1360 7475 1600
rect 8205 1360 8240 1600
rect 7440 980 7475 1220
rect 8205 1050 8240 1290
rect 6845 560 6880 800
rect 7440 510 7475 750
rect 6140 0 6175 240
rect 8205 670 8240 910
rect 8205 395 8240 635
rect 8595 625 8630 865
rect 8595 350 8630 590
rect 8755 625 8790 865
rect 8755 350 8790 590
rect 7440 -10 7475 230
rect 8045 -35 8080 205
rect 8045 -310 8080 -70
rect 8205 -35 8240 205
rect 8205 -310 8240 -70
<< xpolyres >>
rect 5405 240 5440 1360
rect 5565 240 5600 1360
rect 6140 240 6175 1360
rect 6845 800 6880 1360
rect 7440 1220 7475 1360
rect 8205 1290 8240 1360
rect 7440 230 7475 510
rect 8205 635 8240 670
rect 8595 590 8630 625
rect 8755 590 8790 625
rect 8045 -70 8080 -35
rect 8205 -70 8240 -35
<< locali >>
rect 4825 1960 11000 1980
rect 4825 -440 4860 1960
rect 6140 1900 6880 1920
rect 5345 1645 5645 1670
rect 5240 1050 5280 1055
rect 5125 1045 5280 1050
rect 4975 1015 5060 1030
rect 4975 995 4980 1015
rect 5000 995 5020 1015
rect 4975 990 5020 995
rect 5045 990 5060 1015
rect 4975 975 5060 990
rect 5125 1025 5250 1045
rect 5270 1025 5280 1045
rect 4975 930 5000 975
rect 4995 900 5000 930
rect 4975 865 5000 900
rect 4995 835 5000 865
rect 4975 805 5000 835
rect 4995 775 5000 805
rect 4975 740 5000 775
rect 4995 710 5000 740
rect 4975 680 5000 710
rect 4995 650 5000 680
rect 4975 640 5000 650
rect 5025 930 5050 940
rect 5025 900 5030 930
rect 5025 870 5050 900
rect 5025 840 5030 870
rect 5025 805 5050 840
rect 5025 775 5030 805
rect 5025 745 5050 775
rect 5025 715 5030 745
rect 5025 680 5050 715
rect 5025 650 5030 680
rect 5025 615 5050 650
rect 5125 615 5150 1025
rect 5240 1015 5280 1025
rect 5345 995 5370 1645
rect 5440 1360 5565 1600
rect 5180 970 5370 995
rect 5180 835 5205 970
rect 5230 940 5255 950
rect 5250 910 5255 940
rect 5230 890 5255 910
rect 5250 860 5255 890
rect 5230 835 5255 860
rect 5180 810 5255 835
rect 4915 605 4955 615
rect 4915 585 4925 605
rect 4945 585 4955 605
rect 4915 575 4955 585
rect 5025 585 5150 615
rect 5230 780 5255 810
rect 5250 750 5255 780
rect 5230 715 5255 750
rect 5250 685 5255 715
rect 5230 655 5255 685
rect 5250 625 5255 655
rect 5230 590 5255 625
rect 4920 390 4945 575
rect 4975 555 5000 565
rect 4995 525 5000 555
rect 4975 505 5000 525
rect 4995 475 5000 505
rect 4975 445 5000 475
rect 5025 555 5050 585
rect 5025 525 5030 555
rect 5025 505 5050 525
rect 5025 475 5030 505
rect 5250 560 5255 590
rect 5230 530 5255 560
rect 5250 500 5255 530
rect 5230 490 5255 500
rect 5280 940 5305 950
rect 5280 910 5285 940
rect 5280 890 5305 910
rect 5280 860 5285 890
rect 5280 835 5305 860
rect 5280 810 5370 835
rect 5280 780 5305 810
rect 5280 750 5285 780
rect 5280 720 5305 750
rect 5280 690 5285 720
rect 5280 655 5305 690
rect 5280 625 5285 655
rect 5280 595 5305 625
rect 5280 565 5285 595
rect 5280 530 5305 565
rect 5280 500 5285 530
rect 5280 490 5305 500
rect 5025 465 5050 475
rect 4975 440 5010 445
rect 4975 420 4980 440
rect 5005 420 5010 440
rect 4975 410 5010 420
rect 5250 440 5290 450
rect 5250 420 5260 440
rect 5280 420 5290 440
rect 4915 385 4955 390
rect 5250 385 5290 420
rect 4915 380 5290 385
rect 4915 360 4925 380
rect 4945 360 5290 380
rect 4915 355 5290 360
rect 4915 350 4955 355
rect 5345 0 5370 810
rect 5345 -25 5440 0
rect 5405 -440 5440 -25
rect 4825 -470 5440 -440
rect 4830 -475 5440 -470
rect 5620 0 5645 1645
rect 6140 1625 6175 1900
rect 6845 1625 6880 1900
rect 7440 1900 8240 1920
rect 7260 1825 7300 1830
rect 7145 1820 7300 1825
rect 6080 1600 6175 1625
rect 5985 1050 6025 1055
rect 5870 1045 6025 1050
rect 5720 1015 5805 1030
rect 5720 995 5725 1015
rect 5745 995 5765 1015
rect 5720 990 5765 995
rect 5790 990 5805 1015
rect 5720 975 5805 990
rect 5870 1025 5995 1045
rect 6015 1025 6025 1045
rect 5720 930 5745 975
rect 5740 900 5745 930
rect 5720 865 5745 900
rect 5740 835 5745 865
rect 5720 805 5745 835
rect 5740 775 5745 805
rect 5720 740 5745 775
rect 5740 710 5745 740
rect 5720 680 5745 710
rect 5740 650 5745 680
rect 5720 640 5745 650
rect 5770 930 5795 940
rect 5770 900 5775 930
rect 5770 870 5795 900
rect 5770 840 5775 870
rect 5770 805 5795 840
rect 5770 775 5775 805
rect 5770 745 5795 775
rect 5770 715 5775 745
rect 5770 680 5795 715
rect 5770 650 5775 680
rect 5770 615 5795 650
rect 5870 615 5895 1025
rect 5985 1015 6025 1025
rect 6080 995 6105 1600
rect 6720 1600 6880 1625
rect 6590 1050 6630 1055
rect 6475 1045 6630 1050
rect 5925 970 6105 995
rect 6325 1015 6410 1030
rect 6325 995 6330 1015
rect 6350 995 6370 1015
rect 6325 990 6370 995
rect 6395 990 6410 1015
rect 6325 975 6410 990
rect 6475 1025 6600 1045
rect 6620 1025 6630 1045
rect 5925 835 5950 970
rect 5975 940 6000 950
rect 5995 910 6000 940
rect 5975 890 6000 910
rect 5995 860 6000 890
rect 5975 835 6000 860
rect 5925 810 6000 835
rect 5665 605 5705 615
rect 5665 585 5675 605
rect 5695 585 5705 605
rect 5665 575 5705 585
rect 5770 585 5895 615
rect 5975 780 6000 810
rect 5995 750 6000 780
rect 5975 715 6000 750
rect 5995 685 6000 715
rect 5975 655 6000 685
rect 5995 625 6000 655
rect 5975 590 6000 625
rect 5670 390 5695 575
rect 5720 555 5745 565
rect 5740 525 5745 555
rect 5720 505 5745 525
rect 5740 475 5745 505
rect 5720 445 5745 475
rect 5770 555 5795 585
rect 5770 525 5775 555
rect 5770 505 5795 525
rect 5770 475 5775 505
rect 5995 560 6000 590
rect 5975 530 6000 560
rect 5995 500 6000 530
rect 5975 490 6000 500
rect 6025 940 6050 950
rect 6025 910 6030 940
rect 6025 890 6050 910
rect 6025 860 6030 890
rect 6025 835 6050 860
rect 6325 930 6350 975
rect 6345 900 6350 930
rect 6325 865 6350 900
rect 6345 835 6350 865
rect 6025 810 6105 835
rect 6025 780 6050 810
rect 6025 750 6030 780
rect 6025 720 6050 750
rect 6025 690 6030 720
rect 6025 655 6050 690
rect 6025 625 6030 655
rect 6025 595 6050 625
rect 6025 565 6030 595
rect 6025 530 6050 565
rect 6025 500 6030 530
rect 6025 490 6050 500
rect 5770 465 5795 475
rect 5720 440 5755 445
rect 5720 420 5725 440
rect 5750 420 5755 440
rect 5720 410 5755 420
rect 5995 440 6035 450
rect 5995 420 6005 440
rect 6025 420 6035 440
rect 5665 385 5705 390
rect 5995 385 6035 420
rect 5665 380 6035 385
rect 5665 360 5675 380
rect 5695 360 6035 380
rect 5665 355 6035 360
rect 5665 350 5705 355
rect 5565 -25 5645 0
rect 6080 0 6105 810
rect 6325 805 6350 835
rect 6345 775 6350 805
rect 6325 740 6350 775
rect 6345 710 6350 740
rect 6325 680 6350 710
rect 6345 650 6350 680
rect 6325 640 6350 650
rect 6375 930 6400 940
rect 6375 900 6380 930
rect 6375 870 6400 900
rect 6375 840 6380 870
rect 6375 805 6400 840
rect 6375 775 6380 805
rect 6375 745 6400 775
rect 6375 715 6380 745
rect 6375 680 6400 715
rect 6375 650 6380 680
rect 6375 615 6400 650
rect 6475 615 6500 1025
rect 6590 1015 6630 1025
rect 6720 995 6745 1600
rect 6995 1790 7080 1805
rect 6995 1770 7000 1790
rect 7020 1770 7040 1790
rect 6995 1765 7040 1770
rect 7065 1765 7080 1790
rect 6995 1750 7080 1765
rect 7145 1800 7270 1820
rect 7290 1800 7300 1820
rect 6995 1705 7020 1750
rect 7015 1675 7020 1705
rect 6995 1640 7020 1675
rect 7015 1610 7020 1640
rect 6995 1580 7020 1610
rect 7015 1550 7020 1580
rect 6995 1515 7020 1550
rect 7015 1485 7020 1515
rect 6995 1455 7020 1485
rect 7015 1425 7020 1455
rect 6995 1415 7020 1425
rect 7045 1705 7070 1715
rect 7045 1675 7050 1705
rect 7045 1645 7070 1675
rect 7045 1615 7050 1645
rect 7045 1580 7070 1615
rect 7045 1550 7050 1580
rect 7045 1520 7070 1550
rect 7045 1490 7050 1520
rect 7045 1455 7070 1490
rect 7045 1425 7050 1455
rect 7045 1390 7070 1425
rect 7145 1390 7170 1800
rect 7260 1790 7300 1800
rect 7440 1770 7475 1900
rect 7855 1825 7895 1830
rect 7740 1820 7895 1825
rect 7200 1750 7475 1770
rect 7200 1610 7225 1750
rect 7250 1715 7275 1725
rect 7270 1685 7275 1715
rect 7250 1665 7275 1685
rect 7270 1635 7275 1665
rect 7250 1610 7275 1635
rect 7200 1585 7275 1610
rect 6935 1380 6975 1390
rect 6935 1360 6945 1380
rect 6965 1360 6975 1380
rect 6935 1350 6975 1360
rect 7045 1360 7170 1390
rect 7250 1555 7275 1585
rect 7270 1525 7275 1555
rect 7250 1490 7275 1525
rect 7270 1460 7275 1490
rect 7250 1430 7275 1460
rect 7270 1400 7275 1430
rect 7250 1365 7275 1400
rect 6940 1165 6965 1350
rect 6995 1330 7020 1340
rect 7015 1300 7020 1330
rect 6995 1280 7020 1300
rect 7015 1250 7020 1280
rect 6995 1220 7020 1250
rect 7045 1330 7070 1360
rect 7045 1300 7050 1330
rect 7045 1280 7070 1300
rect 7045 1250 7050 1280
rect 7270 1335 7275 1365
rect 7250 1305 7275 1335
rect 7270 1275 7275 1305
rect 7250 1265 7275 1275
rect 7300 1715 7325 1725
rect 7300 1685 7305 1715
rect 7300 1665 7325 1685
rect 7300 1635 7305 1665
rect 7300 1610 7325 1635
rect 7300 1585 7400 1610
rect 7300 1555 7325 1585
rect 7300 1525 7305 1555
rect 7300 1495 7325 1525
rect 7300 1465 7305 1495
rect 7300 1430 7325 1465
rect 7300 1400 7305 1430
rect 7300 1370 7325 1400
rect 7300 1340 7305 1370
rect 7300 1305 7325 1340
rect 7300 1275 7305 1305
rect 7300 1265 7325 1275
rect 7045 1240 7070 1250
rect 6995 1215 7030 1220
rect 6995 1195 7000 1215
rect 7025 1195 7030 1215
rect 6995 1185 7030 1195
rect 7270 1215 7310 1225
rect 7270 1195 7280 1215
rect 7300 1195 7310 1215
rect 6935 1160 6975 1165
rect 7270 1160 7310 1195
rect 6935 1155 7310 1160
rect 6935 1135 6945 1155
rect 6965 1135 7310 1155
rect 6935 1130 7310 1135
rect 6935 1125 6975 1130
rect 7255 1055 7295 1060
rect 7140 1050 7295 1055
rect 6530 970 6745 995
rect 6990 1020 7075 1035
rect 6990 1000 6995 1020
rect 7015 1000 7035 1020
rect 6990 995 7035 1000
rect 7060 995 7075 1020
rect 6990 975 7075 995
rect 7140 1030 7265 1050
rect 7285 1030 7295 1050
rect 6530 835 6555 970
rect 6580 940 6605 950
rect 6600 910 6605 940
rect 6580 890 6605 910
rect 6600 860 6605 890
rect 6580 835 6605 860
rect 6530 810 6605 835
rect 6265 605 6305 615
rect 6265 585 6275 605
rect 6295 585 6305 605
rect 6265 575 6305 585
rect 6375 585 6500 615
rect 6580 780 6605 810
rect 6600 750 6605 780
rect 6580 715 6605 750
rect 6600 685 6605 715
rect 6580 655 6605 685
rect 6600 625 6605 655
rect 6580 590 6605 625
rect 6270 390 6295 575
rect 6325 555 6350 565
rect 6345 525 6350 555
rect 6325 505 6350 525
rect 6345 475 6350 505
rect 6325 445 6350 475
rect 6375 555 6400 585
rect 6375 525 6380 555
rect 6375 505 6400 525
rect 6375 475 6380 505
rect 6600 560 6605 590
rect 6580 530 6605 560
rect 6600 500 6605 530
rect 6580 490 6605 500
rect 6630 940 6655 950
rect 6630 910 6635 940
rect 6630 890 6655 910
rect 6630 860 6635 890
rect 6630 835 6655 860
rect 6990 935 7015 975
rect 7010 905 7015 935
rect 6990 870 7015 905
rect 7010 840 7015 870
rect 6630 810 6715 835
rect 6630 780 6655 810
rect 6630 750 6635 780
rect 6630 720 6655 750
rect 6630 690 6635 720
rect 6630 655 6655 690
rect 6630 625 6635 655
rect 6630 595 6655 625
rect 6630 565 6635 595
rect 6630 530 6655 565
rect 6630 500 6635 530
rect 6690 545 6715 810
rect 6990 810 7015 840
rect 7010 780 7015 810
rect 6990 745 7015 780
rect 7010 715 7015 745
rect 6990 685 7015 715
rect 7010 655 7015 685
rect 6990 645 7015 655
rect 7040 935 7065 945
rect 7040 905 7045 935
rect 7040 875 7065 905
rect 7040 845 7045 875
rect 7040 810 7065 845
rect 7040 780 7045 810
rect 7040 750 7065 780
rect 7040 720 7045 750
rect 7040 685 7065 720
rect 7040 655 7045 685
rect 7040 620 7065 655
rect 7140 620 7165 1030
rect 7255 1020 7295 1030
rect 7375 1000 7400 1585
rect 7440 1600 7475 1750
rect 7590 1790 7675 1805
rect 7590 1770 7595 1790
rect 7615 1770 7635 1790
rect 7590 1765 7635 1770
rect 7660 1765 7675 1790
rect 7590 1750 7675 1765
rect 7740 1800 7865 1820
rect 7885 1800 7895 1820
rect 7590 1705 7615 1750
rect 7610 1675 7615 1705
rect 7590 1640 7615 1675
rect 7610 1610 7615 1640
rect 7590 1580 7615 1610
rect 7610 1550 7615 1580
rect 7590 1515 7615 1550
rect 7610 1485 7615 1515
rect 7590 1455 7615 1485
rect 7610 1425 7615 1455
rect 7590 1415 7615 1425
rect 7640 1705 7665 1715
rect 7640 1675 7645 1705
rect 7640 1645 7665 1675
rect 7640 1615 7645 1645
rect 7640 1580 7665 1615
rect 7640 1550 7645 1580
rect 7640 1520 7665 1550
rect 7640 1490 7645 1520
rect 7640 1455 7665 1490
rect 7640 1425 7645 1455
rect 7640 1390 7665 1425
rect 7740 1390 7765 1800
rect 7855 1790 7895 1800
rect 8205 1770 8240 1900
rect 8620 1900 8755 1915
rect 8620 1865 8635 1900
rect 8660 1865 8720 1900
rect 8745 1865 8755 1900
rect 8620 1855 8755 1865
rect 8895 1900 8985 1915
rect 8895 1865 8905 1900
rect 8930 1865 8950 1900
rect 8975 1865 8985 1900
rect 7795 1750 8240 1770
rect 7795 1610 7820 1750
rect 7845 1715 7870 1725
rect 7865 1685 7870 1715
rect 7845 1665 7870 1685
rect 7865 1635 7870 1665
rect 7845 1610 7870 1635
rect 7795 1585 7870 1610
rect 7530 1380 7570 1390
rect 7530 1360 7540 1380
rect 7560 1360 7570 1380
rect 7530 1350 7570 1360
rect 7640 1360 7765 1390
rect 7845 1555 7870 1585
rect 7865 1525 7870 1555
rect 7845 1490 7870 1525
rect 7865 1460 7870 1490
rect 7845 1430 7870 1460
rect 7865 1400 7870 1430
rect 7845 1365 7870 1400
rect 7195 975 7400 1000
rect 7535 1165 7560 1350
rect 7590 1330 7615 1340
rect 7610 1300 7615 1330
rect 7590 1280 7615 1300
rect 7610 1250 7615 1280
rect 7590 1220 7615 1250
rect 7640 1330 7665 1360
rect 7640 1300 7645 1330
rect 7640 1280 7665 1300
rect 7640 1250 7645 1280
rect 7865 1335 7870 1365
rect 7845 1305 7870 1335
rect 7865 1275 7870 1305
rect 7845 1265 7870 1275
rect 7895 1715 7920 1725
rect 7895 1685 7900 1715
rect 7895 1665 7920 1685
rect 7895 1635 7900 1665
rect 7895 1610 7920 1635
rect 7895 1585 7995 1610
rect 7895 1555 7920 1585
rect 7895 1525 7900 1555
rect 7895 1495 7920 1525
rect 7895 1465 7900 1495
rect 7895 1430 7920 1465
rect 7895 1400 7900 1430
rect 7895 1370 7920 1400
rect 7895 1340 7900 1370
rect 7895 1305 7920 1340
rect 7895 1275 7900 1305
rect 7895 1265 7920 1275
rect 7640 1240 7665 1250
rect 7590 1215 7625 1220
rect 7590 1195 7595 1215
rect 7620 1195 7625 1215
rect 7590 1185 7625 1195
rect 7865 1215 7905 1225
rect 7865 1195 7875 1215
rect 7895 1195 7905 1215
rect 7530 1160 7570 1165
rect 7865 1160 7905 1195
rect 7530 1155 7905 1160
rect 7530 1135 7540 1155
rect 7560 1135 7905 1155
rect 7530 1130 7905 1135
rect 7530 1125 7570 1130
rect 7850 1055 7890 1060
rect 7735 1050 7890 1055
rect 7440 975 7475 980
rect 7195 840 7220 975
rect 7245 945 7270 955
rect 7265 915 7270 945
rect 7245 895 7270 915
rect 7265 865 7270 895
rect 7245 840 7270 865
rect 7195 815 7270 840
rect 6930 610 6970 620
rect 6930 590 6940 610
rect 6960 590 6970 610
rect 6930 580 6970 590
rect 7040 590 7165 620
rect 7245 785 7270 815
rect 7265 755 7270 785
rect 7245 720 7270 755
rect 7265 690 7270 720
rect 7245 660 7270 690
rect 7265 630 7270 660
rect 7245 595 7270 630
rect 6845 545 6880 560
rect 6690 520 6880 545
rect 6630 490 6655 500
rect 6375 465 6400 475
rect 6325 440 6360 445
rect 6325 420 6330 440
rect 6355 420 6360 440
rect 6325 410 6360 420
rect 6600 440 6640 450
rect 6600 420 6610 440
rect 6630 420 6640 440
rect 6265 385 6305 390
rect 6600 385 6640 420
rect 6265 380 6640 385
rect 6265 360 6275 380
rect 6295 360 6640 380
rect 6265 355 6640 360
rect 6265 350 6305 355
rect 6080 -25 6175 0
rect 5565 -520 5600 -25
rect 6140 -520 6175 -25
rect 5565 -555 6175 -520
rect 6845 -520 6880 520
rect 6935 395 6960 580
rect 6990 560 7015 570
rect 7010 530 7015 560
rect 6990 510 7015 530
rect 7010 480 7015 510
rect 6990 450 7015 480
rect 7040 560 7065 590
rect 7040 530 7045 560
rect 7040 510 7065 530
rect 7040 480 7045 510
rect 7265 565 7270 595
rect 7245 535 7270 565
rect 7265 505 7270 535
rect 7245 495 7270 505
rect 7295 945 7320 955
rect 7375 950 7475 975
rect 7295 915 7300 945
rect 7295 895 7320 915
rect 7295 865 7300 895
rect 7295 840 7320 865
rect 7295 815 7395 840
rect 7295 785 7320 815
rect 7295 755 7300 785
rect 7295 725 7320 755
rect 7295 695 7300 725
rect 7295 660 7320 695
rect 7295 630 7300 660
rect 7295 600 7320 630
rect 7295 570 7300 600
rect 7295 535 7320 570
rect 7295 505 7300 535
rect 7295 495 7320 505
rect 7040 470 7065 480
rect 6990 445 7025 450
rect 6990 425 6995 445
rect 7020 425 7025 445
rect 6990 415 7025 425
rect 7265 445 7305 455
rect 7265 425 7275 445
rect 7295 425 7305 445
rect 6930 390 6970 395
rect 7265 390 7305 425
rect 6930 385 7305 390
rect 6930 365 6940 385
rect 6960 365 7305 385
rect 6930 360 7305 365
rect 6930 355 6970 360
rect 7370 -25 7395 815
rect 7440 750 7475 950
rect 7585 1020 7670 1035
rect 7585 1000 7590 1020
rect 7610 1000 7630 1020
rect 7585 995 7630 1000
rect 7655 995 7670 1020
rect 7585 980 7670 995
rect 7735 1030 7860 1050
rect 7880 1030 7890 1050
rect 7585 935 7610 980
rect 7605 905 7610 935
rect 7585 870 7610 905
rect 7605 840 7610 870
rect 7585 810 7610 840
rect 7605 780 7610 810
rect 7585 745 7610 780
rect 7605 715 7610 745
rect 7585 685 7610 715
rect 7605 655 7610 685
rect 7585 645 7610 655
rect 7635 935 7660 945
rect 7635 905 7640 935
rect 7635 875 7660 905
rect 7635 845 7640 875
rect 7635 810 7660 845
rect 7635 780 7640 810
rect 7635 750 7660 780
rect 7635 720 7640 750
rect 7635 685 7660 720
rect 7635 655 7640 685
rect 7635 620 7660 655
rect 7735 620 7760 1030
rect 7850 1020 7890 1030
rect 7970 1000 7995 1585
rect 8205 1600 8240 1750
rect 8205 1000 8240 1050
rect 7790 975 8240 1000
rect 7790 840 7815 975
rect 7840 945 7865 955
rect 7860 915 7865 945
rect 7840 895 7865 915
rect 7860 865 7865 895
rect 7840 840 7865 865
rect 7790 815 7865 840
rect 7525 610 7565 620
rect 7525 590 7535 610
rect 7555 590 7565 610
rect 7525 580 7565 590
rect 7635 590 7760 620
rect 7840 785 7865 815
rect 7860 755 7865 785
rect 7840 720 7865 755
rect 7860 690 7865 720
rect 7840 660 7865 690
rect 7860 630 7865 660
rect 7840 595 7865 630
rect 7530 395 7555 580
rect 7585 560 7610 570
rect 7605 530 7610 560
rect 7585 510 7610 530
rect 7605 480 7610 510
rect 7585 450 7610 480
rect 7635 560 7660 590
rect 7635 530 7640 560
rect 7635 510 7660 530
rect 7635 480 7640 510
rect 7860 565 7865 595
rect 7840 535 7865 565
rect 7860 505 7865 535
rect 7840 495 7865 505
rect 7890 945 7915 955
rect 7890 915 7895 945
rect 7890 895 7915 915
rect 7890 865 7895 895
rect 7890 840 7915 865
rect 8205 910 8240 975
rect 7890 815 7990 840
rect 7890 785 7915 815
rect 7890 755 7895 785
rect 7890 725 7915 755
rect 7890 695 7895 725
rect 7890 660 7915 695
rect 7890 630 7895 660
rect 7890 600 7915 630
rect 7890 570 7895 600
rect 7890 535 7915 570
rect 7890 505 7895 535
rect 7890 495 7915 505
rect 7635 470 7660 480
rect 7585 445 7620 450
rect 7585 425 7590 445
rect 7615 425 7620 445
rect 7585 415 7620 425
rect 7860 445 7900 455
rect 7860 425 7870 445
rect 7890 425 7900 445
rect 7525 390 7565 395
rect 7860 390 7900 425
rect 7525 385 7900 390
rect 7525 365 7535 385
rect 7555 365 7900 385
rect 7525 360 7900 365
rect 7525 355 7565 360
rect 7965 295 7990 815
rect 8665 865 8715 1855
rect 8895 1600 8985 1865
rect 9500 1750 10680 1780
rect 9540 1710 9560 1750
rect 9600 1710 9620 1750
rect 9660 1710 9680 1750
rect 9720 1710 9740 1750
rect 9780 1710 9800 1750
rect 9840 1710 9860 1750
rect 9900 1710 9920 1750
rect 9960 1710 9980 1750
rect 10020 1710 10040 1750
rect 10080 1710 10100 1750
rect 10140 1710 10160 1750
rect 10200 1710 10220 1750
rect 10260 1710 10280 1750
rect 10320 1710 10340 1750
rect 10380 1710 10400 1750
rect 10440 1710 10460 1750
rect 10500 1710 10520 1750
rect 10560 1730 10680 1750
rect 10560 1710 10600 1730
rect 9500 1690 10600 1710
rect 9540 1650 9560 1690
rect 9600 1650 9620 1690
rect 9660 1650 9680 1690
rect 9720 1650 9740 1690
rect 9780 1650 9800 1690
rect 9840 1650 9860 1690
rect 9900 1650 9920 1690
rect 9960 1650 9980 1690
rect 10020 1650 10040 1690
rect 10080 1650 10100 1690
rect 10140 1650 10160 1690
rect 10200 1650 10220 1690
rect 10260 1650 10280 1690
rect 10320 1650 10340 1690
rect 10380 1650 10400 1690
rect 10440 1650 10460 1690
rect 10500 1650 10520 1690
rect 10560 1670 10600 1690
rect 10650 1670 10680 1730
rect 10560 1650 10680 1670
rect 9500 1620 10680 1650
rect 8895 1565 8905 1600
rect 8930 1565 8950 1600
rect 8975 1565 8985 1600
rect 8895 1555 8985 1565
rect 9370 1510 9420 1560
rect 9370 1480 9380 1510
rect 9410 1480 9420 1510
rect 9370 1460 9420 1480
rect 9370 1430 9380 1460
rect 9410 1430 9420 1460
rect 9370 1410 9420 1430
rect 9370 1380 9380 1410
rect 9410 1380 9420 1410
rect 9370 1360 9420 1380
rect 9370 1330 9380 1360
rect 9410 1330 9420 1360
rect 9370 1310 9420 1330
rect 9370 1280 9380 1310
rect 9410 1280 9420 1310
rect 9370 1260 9420 1280
rect 9370 1230 9380 1260
rect 9410 1230 9420 1260
rect 9370 1210 9420 1230
rect 9370 1180 9380 1210
rect 9410 1180 9420 1210
rect 9370 1160 9420 1180
rect 9370 1130 9380 1160
rect 9410 1130 9420 1160
rect 9370 1110 9420 1130
rect 9370 1080 9380 1110
rect 9410 1080 9420 1110
rect 9370 1060 9420 1080
rect 9370 1030 9380 1060
rect 9410 1030 9420 1060
rect 9370 1010 9420 1030
rect 9370 980 9380 1010
rect 9410 980 9420 1010
rect 9370 920 9420 980
rect 9520 1510 9570 1620
rect 9520 1480 9530 1510
rect 9560 1480 9570 1510
rect 9520 1460 9570 1480
rect 9520 1430 9530 1460
rect 9560 1430 9570 1460
rect 9520 1410 9570 1430
rect 9520 1380 9530 1410
rect 9560 1380 9570 1410
rect 9520 1360 9570 1380
rect 9520 1330 9530 1360
rect 9560 1330 9570 1360
rect 9520 1310 9570 1330
rect 9520 1280 9530 1310
rect 9560 1280 9570 1310
rect 9520 1260 9570 1280
rect 9520 1230 9530 1260
rect 9560 1230 9570 1260
rect 9520 1210 9570 1230
rect 9520 1180 9530 1210
rect 9560 1180 9570 1210
rect 9520 1160 9570 1180
rect 9520 1130 9530 1160
rect 9560 1130 9570 1160
rect 9520 1110 9570 1130
rect 9520 1080 9530 1110
rect 9560 1080 9570 1110
rect 9520 1060 9570 1080
rect 9520 1030 9530 1060
rect 9560 1030 9570 1060
rect 9520 1010 9570 1030
rect 9520 980 9530 1010
rect 9560 980 9570 1010
rect 9520 940 9570 980
rect 9670 1510 9720 1560
rect 9670 1480 9680 1510
rect 9710 1480 9720 1510
rect 9670 1460 9720 1480
rect 9670 1430 9680 1460
rect 9710 1430 9720 1460
rect 9670 1410 9720 1430
rect 9670 1380 9680 1410
rect 9710 1380 9720 1410
rect 9670 1360 9720 1380
rect 9670 1330 9680 1360
rect 9710 1330 9720 1360
rect 9670 1310 9720 1330
rect 9670 1280 9680 1310
rect 9710 1280 9720 1310
rect 9670 1260 9720 1280
rect 9670 1230 9680 1260
rect 9710 1230 9720 1260
rect 9670 1210 9720 1230
rect 9670 1180 9680 1210
rect 9710 1180 9720 1210
rect 9670 1160 9720 1180
rect 9670 1130 9680 1160
rect 9710 1130 9720 1160
rect 9670 1110 9720 1130
rect 9670 1080 9680 1110
rect 9710 1080 9720 1110
rect 9670 1060 9720 1080
rect 9670 1030 9680 1060
rect 9710 1030 9720 1060
rect 9670 1010 9720 1030
rect 9670 980 9680 1010
rect 9710 980 9720 1010
rect 9370 910 9470 920
rect 9370 870 9430 910
rect 9460 870 9470 910
rect 8630 625 8755 865
rect 9370 860 9470 870
rect 9060 830 9170 850
rect 9420 830 9470 860
rect 9060 770 9470 830
rect 9670 820 9720 980
rect 9770 1510 9820 1560
rect 9770 1480 9780 1510
rect 9810 1480 9820 1510
rect 9770 1460 9820 1480
rect 9770 1430 9780 1460
rect 9810 1430 9820 1460
rect 9770 1410 9820 1430
rect 9770 1380 9780 1410
rect 9810 1380 9820 1410
rect 9770 1360 9820 1380
rect 9770 1330 9780 1360
rect 9810 1330 9820 1360
rect 9770 1310 9820 1330
rect 9770 1280 9780 1310
rect 9810 1280 9820 1310
rect 9770 1260 9820 1280
rect 9770 1230 9780 1260
rect 9810 1230 9820 1260
rect 9770 1210 9820 1230
rect 9770 1180 9780 1210
rect 9810 1180 9820 1210
rect 9770 1160 9820 1180
rect 9770 1130 9780 1160
rect 9810 1130 9820 1160
rect 9770 1110 9820 1130
rect 9770 1080 9780 1110
rect 9810 1080 9820 1110
rect 9770 1060 9820 1080
rect 9770 1030 9780 1060
rect 9810 1030 9820 1060
rect 9770 1010 9820 1030
rect 9770 980 9780 1010
rect 9810 980 9820 1010
rect 9770 910 9820 980
rect 9920 1510 9970 1620
rect 9920 1480 9930 1510
rect 9960 1480 9970 1510
rect 9920 1460 9970 1480
rect 9920 1430 9930 1460
rect 9960 1430 9970 1460
rect 9920 1410 9970 1430
rect 9920 1380 9930 1410
rect 9960 1380 9970 1410
rect 9920 1360 9970 1380
rect 9920 1330 9930 1360
rect 9960 1330 9970 1360
rect 9920 1310 9970 1330
rect 9920 1280 9930 1310
rect 9960 1280 9970 1310
rect 9920 1260 9970 1280
rect 9920 1230 9930 1260
rect 9960 1230 9970 1260
rect 9920 1210 9970 1230
rect 9920 1180 9930 1210
rect 9960 1180 9970 1210
rect 9920 1160 9970 1180
rect 9920 1130 9930 1160
rect 9960 1130 9970 1160
rect 9920 1110 9970 1130
rect 9920 1080 9930 1110
rect 9960 1080 9970 1110
rect 9920 1060 9970 1080
rect 9920 1030 9930 1060
rect 9960 1030 9970 1060
rect 9920 1010 9970 1030
rect 9920 980 9930 1010
rect 9960 980 9970 1010
rect 9920 940 9970 980
rect 10070 1510 10120 1560
rect 10070 1480 10080 1510
rect 10110 1480 10120 1510
rect 10070 1460 10120 1480
rect 10070 1430 10080 1460
rect 10110 1430 10120 1460
rect 10070 1410 10120 1430
rect 10070 1380 10080 1410
rect 10110 1380 10120 1410
rect 10070 1360 10120 1380
rect 10070 1330 10080 1360
rect 10110 1330 10120 1360
rect 10070 1310 10120 1330
rect 10070 1280 10080 1310
rect 10110 1280 10120 1310
rect 10070 1260 10120 1280
rect 10070 1230 10080 1260
rect 10110 1230 10120 1260
rect 10070 1210 10120 1230
rect 10070 1180 10080 1210
rect 10110 1180 10120 1210
rect 10070 1160 10120 1180
rect 10070 1130 10080 1160
rect 10110 1130 10120 1160
rect 10070 1110 10120 1130
rect 10070 1080 10080 1110
rect 10110 1080 10120 1110
rect 10070 1060 10120 1080
rect 10070 1030 10080 1060
rect 10110 1030 10120 1060
rect 10070 1010 10120 1030
rect 10070 980 10080 1010
rect 10110 980 10120 1010
rect 10070 910 10120 980
rect 10220 1510 10270 1620
rect 10220 1480 10230 1510
rect 10260 1480 10270 1510
rect 10220 1460 10270 1480
rect 10220 1430 10230 1460
rect 10260 1430 10270 1460
rect 10220 1410 10270 1430
rect 10220 1380 10230 1410
rect 10260 1380 10270 1410
rect 10220 1360 10270 1380
rect 10220 1330 10230 1360
rect 10260 1330 10270 1360
rect 10220 1310 10270 1330
rect 10220 1280 10230 1310
rect 10260 1280 10270 1310
rect 10220 1260 10270 1280
rect 10220 1230 10230 1260
rect 10260 1230 10270 1260
rect 10220 1210 10270 1230
rect 10220 1180 10230 1210
rect 10260 1180 10270 1210
rect 10220 1160 10270 1180
rect 10220 1130 10230 1160
rect 10260 1130 10270 1160
rect 10220 1110 10270 1130
rect 10220 1080 10230 1110
rect 10260 1080 10270 1110
rect 10220 1060 10270 1080
rect 10220 1030 10230 1060
rect 10260 1030 10270 1060
rect 10220 1010 10270 1030
rect 10220 980 10230 1010
rect 10260 980 10270 1010
rect 10220 940 10270 980
rect 10370 1510 10420 1560
rect 10370 1480 10380 1510
rect 10410 1480 10420 1510
rect 10370 1460 10420 1480
rect 10370 1430 10380 1460
rect 10410 1430 10420 1460
rect 10370 1410 10420 1430
rect 10370 1380 10380 1410
rect 10410 1380 10420 1410
rect 10370 1360 10420 1380
rect 10370 1330 10380 1360
rect 10410 1330 10420 1360
rect 10370 1310 10420 1330
rect 10370 1280 10380 1310
rect 10410 1280 10420 1310
rect 10370 1260 10420 1280
rect 10370 1230 10380 1260
rect 10410 1230 10420 1260
rect 10370 1210 10420 1230
rect 10370 1180 10380 1210
rect 10410 1180 10420 1210
rect 10370 1160 10420 1180
rect 10370 1130 10380 1160
rect 10410 1130 10420 1160
rect 10370 1110 10420 1130
rect 10370 1080 10380 1110
rect 10410 1080 10420 1110
rect 10370 1060 10420 1080
rect 10370 1030 10380 1060
rect 10410 1030 10420 1060
rect 10370 1010 10420 1030
rect 10370 980 10380 1010
rect 10410 980 10420 1010
rect 10370 910 10420 980
rect 10520 1510 10570 1620
rect 10520 1480 10530 1510
rect 10560 1480 10570 1510
rect 10520 1460 10570 1480
rect 10520 1430 10530 1460
rect 10560 1430 10570 1460
rect 10520 1410 10570 1430
rect 10520 1380 10530 1410
rect 10560 1380 10570 1410
rect 10520 1360 10570 1380
rect 10520 1330 10530 1360
rect 10560 1330 10570 1360
rect 10520 1310 10570 1330
rect 10520 1280 10530 1310
rect 10560 1280 10570 1310
rect 10520 1260 10570 1280
rect 10520 1230 10530 1260
rect 10560 1230 10570 1260
rect 10520 1210 10570 1230
rect 10520 1180 10530 1210
rect 10560 1180 10570 1210
rect 10520 1160 10570 1180
rect 10520 1130 10530 1160
rect 10560 1130 10570 1160
rect 10520 1110 10570 1130
rect 10520 1080 10530 1110
rect 10560 1080 10570 1110
rect 10520 1060 10570 1080
rect 10520 1030 10530 1060
rect 10560 1030 10570 1060
rect 10520 1010 10570 1030
rect 10520 980 10530 1010
rect 10560 980 10570 1010
rect 10520 940 10570 980
rect 10670 1510 10720 1560
rect 10670 1480 10680 1510
rect 10710 1480 10720 1510
rect 10670 1460 10720 1480
rect 10670 1430 10680 1460
rect 10710 1430 10720 1460
rect 10670 1410 10720 1430
rect 10670 1380 10680 1410
rect 10710 1380 10720 1410
rect 10670 1360 10720 1380
rect 10670 1330 10680 1360
rect 10710 1330 10720 1360
rect 10670 1310 10720 1330
rect 10670 1280 10680 1310
rect 10710 1280 10720 1310
rect 10670 1260 10720 1280
rect 10670 1230 10680 1260
rect 10710 1230 10720 1260
rect 10670 1210 10720 1230
rect 10670 1180 10680 1210
rect 10710 1180 10720 1210
rect 10670 1160 10720 1180
rect 10670 1130 10680 1160
rect 10710 1130 10720 1160
rect 10670 1110 10720 1130
rect 10670 1080 10680 1110
rect 10710 1080 10720 1110
rect 10670 1060 10720 1080
rect 10670 1030 10680 1060
rect 10710 1030 10720 1060
rect 10670 1010 10720 1030
rect 10670 980 10680 1010
rect 10710 980 10720 1010
rect 9770 860 10420 910
rect 9520 770 9720 820
rect 10110 795 10220 810
rect 9060 750 9170 770
rect 9370 660 9420 680
rect 9370 630 9380 660
rect 9410 630 9420 660
rect 9370 610 9420 630
rect 8205 295 8240 395
rect 7965 270 8240 295
rect 8630 330 8755 590
rect 9370 580 9380 610
rect 9410 580 9420 610
rect 9370 560 9420 580
rect 9370 530 9380 560
rect 9410 530 9420 560
rect 9370 510 9420 530
rect 9370 480 9380 510
rect 9410 480 9420 510
rect 9370 460 9420 480
rect 9370 400 9380 460
rect 9410 400 9420 460
rect 9030 340 9140 350
rect 9030 330 9040 340
rect 8630 270 9040 330
rect 7850 245 7890 250
rect 7735 240 7890 245
rect 7440 -25 7475 -10
rect 7370 -50 7475 -25
rect 7440 -520 7475 -50
rect 7585 210 7670 225
rect 7585 190 7590 210
rect 7610 190 7630 210
rect 7585 185 7630 190
rect 7655 185 7670 210
rect 7585 170 7670 185
rect 7735 220 7860 240
rect 7880 220 7890 240
rect 7585 125 7610 170
rect 7605 95 7610 125
rect 7585 60 7610 95
rect 7605 30 7610 60
rect 7585 0 7610 30
rect 7605 -30 7610 0
rect 7585 -65 7610 -30
rect 7605 -95 7610 -65
rect 7585 -125 7610 -95
rect 7605 -155 7610 -125
rect 7585 -165 7610 -155
rect 7635 125 7660 135
rect 7635 95 7640 125
rect 7635 65 7660 95
rect 7635 35 7640 65
rect 7635 0 7660 35
rect 7635 -30 7640 0
rect 7635 -60 7660 -30
rect 7635 -90 7640 -60
rect 7635 -125 7660 -90
rect 7635 -155 7640 -125
rect 7635 -190 7660 -155
rect 7735 -190 7760 220
rect 7850 210 7890 220
rect 7965 190 7990 270
rect 8205 205 8240 270
rect 7790 165 7990 190
rect 7790 30 7815 165
rect 7840 135 7865 145
rect 7860 105 7865 135
rect 7840 85 7865 105
rect 7860 55 7865 85
rect 7840 30 7865 55
rect 7790 5 7865 30
rect 7525 -200 7565 -190
rect 7525 -220 7535 -200
rect 7555 -220 7565 -200
rect 7525 -230 7565 -220
rect 7635 -220 7760 -190
rect 7840 -25 7865 5
rect 7860 -55 7865 -25
rect 7840 -90 7865 -55
rect 7860 -120 7865 -90
rect 7840 -150 7865 -120
rect 7860 -180 7865 -150
rect 7840 -215 7865 -180
rect 7530 -415 7555 -230
rect 7585 -250 7610 -240
rect 7605 -280 7610 -250
rect 7585 -300 7610 -280
rect 7605 -330 7610 -300
rect 7585 -360 7610 -330
rect 7635 -250 7660 -220
rect 7635 -280 7640 -250
rect 7635 -300 7660 -280
rect 7635 -330 7640 -300
rect 7860 -245 7865 -215
rect 7840 -275 7865 -245
rect 7860 -305 7865 -275
rect 7840 -315 7865 -305
rect 7890 135 7915 145
rect 7890 105 7895 135
rect 7890 85 7915 105
rect 7890 55 7895 85
rect 7890 30 7915 55
rect 7890 5 7990 30
rect 7890 -25 7915 5
rect 7890 -55 7895 -25
rect 7890 -85 7915 -55
rect 7890 -115 7895 -85
rect 7890 -150 7915 -115
rect 7890 -180 7895 -150
rect 7890 -210 7915 -180
rect 7890 -240 7895 -210
rect 7890 -275 7915 -240
rect 7890 -305 7895 -275
rect 7890 -315 7915 -305
rect 7635 -340 7660 -330
rect 7585 -365 7620 -360
rect 7585 -385 7590 -365
rect 7615 -385 7620 -365
rect 7585 -395 7620 -385
rect 7860 -365 7900 -355
rect 7860 -385 7870 -365
rect 7890 -385 7900 -365
rect 7965 -360 7990 5
rect 8080 -35 8205 205
rect 8680 15 8720 270
rect 9030 260 9040 270
rect 9130 260 9140 340
rect 9030 250 9140 260
rect 9030 205 9140 220
rect 9030 130 9040 205
rect 9135 130 9140 205
rect 9030 120 9140 130
rect 8390 -20 8720 15
rect 9370 90 9420 400
rect 9520 660 9570 770
rect 10110 730 10130 795
rect 10195 730 10220 795
rect 10110 710 10220 730
rect 9520 630 9530 660
rect 9560 630 9570 660
rect 9520 610 9570 630
rect 9520 580 9530 610
rect 9560 580 9570 610
rect 9520 560 9570 580
rect 9520 530 9530 560
rect 9560 530 9570 560
rect 9520 510 9570 530
rect 9520 480 9530 510
rect 9560 480 9570 510
rect 9520 460 9570 480
rect 9520 400 9530 460
rect 9560 400 9570 460
rect 9520 380 9570 400
rect 9670 660 9720 680
rect 9670 630 9680 660
rect 9710 630 9720 660
rect 9670 610 9720 630
rect 9670 580 9680 610
rect 9710 580 9720 610
rect 9670 560 9720 580
rect 9670 530 9680 560
rect 9710 530 9720 560
rect 9670 510 9720 530
rect 9670 480 9680 510
rect 9710 480 9720 510
rect 9670 460 9720 480
rect 9670 400 9680 460
rect 9710 400 9720 460
rect 9670 270 9720 400
rect 10140 630 10190 710
rect 10140 600 10150 630
rect 10180 600 10190 630
rect 10140 580 10190 600
rect 10140 550 10150 580
rect 10180 550 10190 580
rect 10140 530 10190 550
rect 10140 500 10150 530
rect 10180 500 10190 530
rect 10140 480 10190 500
rect 10140 450 10150 480
rect 10180 450 10190 480
rect 10140 430 10190 450
rect 10140 400 10150 430
rect 10180 400 10190 430
rect 10140 380 10190 400
rect 10140 350 10150 380
rect 10180 350 10190 380
rect 10140 330 10190 350
rect 10140 300 10150 330
rect 10180 300 10190 330
rect 10140 280 10190 300
rect 9670 220 9940 270
rect 9370 80 9500 90
rect 9370 40 9430 80
rect 9490 40 9500 80
rect 9370 30 9500 40
rect 9370 0 9420 30
rect 8080 -310 8205 -70
rect 8120 -360 8170 -310
rect 7965 -385 8170 -360
rect 7525 -420 7565 -415
rect 7860 -420 7900 -385
rect 7525 -425 7900 -420
rect 7525 -445 7535 -425
rect 7555 -445 7900 -425
rect 8120 -400 8170 -385
rect 8390 -400 8425 -20
rect 9370 -50 9380 0
rect 9410 -50 9420 0
rect 9370 -80 9420 -50
rect 9520 0 9570 10
rect 9520 -50 9530 0
rect 9560 -50 9570 0
rect 9520 -340 9570 -50
rect 9670 0 9720 220
rect 9670 -50 9680 0
rect 9710 -50 9720 0
rect 9670 -80 9720 -50
rect 9890 -230 9940 220
rect 10140 250 10150 280
rect 10180 250 10190 280
rect 10140 230 10190 250
rect 10140 200 10150 230
rect 10180 200 10190 230
rect 10140 180 10190 200
rect 10140 150 10150 180
rect 10180 150 10190 180
rect 10140 130 10190 150
rect 10140 100 10150 130
rect 10180 100 10190 130
rect 10140 80 10190 100
rect 10140 50 10150 80
rect 10180 50 10190 80
rect 10140 30 10190 50
rect 10140 0 10150 30
rect 10180 0 10190 30
rect 10140 -20 10190 0
rect 10140 -50 10150 -20
rect 10180 -50 10190 -20
rect 10140 -70 10190 -50
rect 10140 -100 10150 -70
rect 10180 -100 10190 -70
rect 10140 -120 10190 -100
rect 10140 -150 10150 -120
rect 10180 -150 10190 -120
rect 10140 -170 10190 -150
rect 10140 -200 10150 -170
rect 10180 -200 10190 -170
rect 10140 -210 10190 -200
rect 10290 630 10340 860
rect 10670 800 10720 980
rect 10965 800 11000 1960
rect 11025 800 11130 825
rect 10670 750 11130 800
rect 10290 600 10300 630
rect 10330 600 10340 630
rect 10290 580 10340 600
rect 10290 550 10300 580
rect 10330 550 10340 580
rect 10290 530 10340 550
rect 10290 500 10300 530
rect 10330 500 10340 530
rect 10290 480 10340 500
rect 10290 450 10300 480
rect 10330 450 10340 480
rect 10290 430 10340 450
rect 10290 400 10300 430
rect 10330 400 10340 430
rect 10290 380 10340 400
rect 10290 350 10300 380
rect 10330 350 10340 380
rect 10290 330 10340 350
rect 10290 300 10300 330
rect 10330 300 10340 330
rect 10290 280 10340 300
rect 10290 250 10300 280
rect 10330 250 10340 280
rect 10290 230 10340 250
rect 10290 200 10300 230
rect 10330 200 10340 230
rect 10290 180 10340 200
rect 10290 150 10300 180
rect 10330 150 10340 180
rect 10290 130 10340 150
rect 10290 100 10300 130
rect 10330 100 10340 130
rect 10290 80 10340 100
rect 10290 50 10300 80
rect 10330 50 10340 80
rect 10290 30 10340 50
rect 10720 590 10770 750
rect 11025 725 11130 750
rect 10720 560 10730 590
rect 10760 560 10770 590
rect 10720 540 10770 560
rect 10720 510 10730 540
rect 10760 510 10770 540
rect 10720 490 10770 510
rect 10720 460 10730 490
rect 10760 460 10770 490
rect 10720 440 10770 460
rect 10720 410 10730 440
rect 10760 410 10770 440
rect 10720 390 10770 410
rect 10720 360 10730 390
rect 10760 360 10770 390
rect 10720 340 10770 360
rect 10720 310 10730 340
rect 10760 310 10770 340
rect 10720 290 10770 310
rect 10720 260 10730 290
rect 10760 260 10770 290
rect 10720 240 10770 260
rect 10720 210 10730 240
rect 10760 210 10770 240
rect 10720 190 10770 210
rect 10720 160 10730 190
rect 10760 160 10770 190
rect 10720 140 10770 160
rect 10720 110 10730 140
rect 10760 110 10770 140
rect 10720 90 10770 110
rect 10720 60 10730 90
rect 10760 60 10770 90
rect 10720 41 10770 60
rect 10870 590 10920 621
rect 10870 560 10880 590
rect 10910 560 10920 590
rect 10870 540 10920 560
rect 10870 510 10880 540
rect 10910 510 10920 540
rect 10870 490 10920 510
rect 10870 460 10880 490
rect 10910 460 10920 490
rect 10870 440 10920 460
rect 10870 410 10880 440
rect 10910 410 10920 440
rect 10870 390 10920 410
rect 10870 360 10880 390
rect 10910 360 10920 390
rect 10870 340 10920 360
rect 10870 310 10880 340
rect 10910 310 10920 340
rect 10870 290 10920 310
rect 10870 260 10880 290
rect 10910 260 10920 290
rect 10870 240 10920 260
rect 10870 210 10880 240
rect 10910 210 10920 240
rect 10870 190 10920 210
rect 10870 160 10880 190
rect 10910 160 10920 190
rect 10870 140 10920 160
rect 10870 110 10880 140
rect 10910 110 10920 140
rect 10870 90 10920 110
rect 10870 60 10880 90
rect 10910 60 10920 90
rect 10290 0 10300 30
rect 10330 0 10340 30
rect 10290 -20 10340 0
rect 10290 -50 10300 -20
rect 10330 -50 10340 -20
rect 10290 -70 10340 -50
rect 10290 -100 10300 -70
rect 10330 -100 10340 -70
rect 10290 -120 10340 -100
rect 10290 -150 10300 -120
rect 10330 -150 10340 -120
rect 10290 -170 10340 -150
rect 10290 -200 10300 -170
rect 10330 -200 10340 -170
rect 10290 -230 10340 -200
rect 10770 10 10850 21
rect 10770 -30 10780 10
rect 10840 -30 10850 10
rect 10770 -230 10850 -30
rect 9890 -240 10270 -230
rect 9890 -280 10210 -240
rect 10250 -280 10270 -240
rect 9890 -290 10270 -280
rect 10290 -280 10850 -230
rect 10870 -180 10920 60
rect 10870 -200 11045 -180
rect 10870 -260 10890 -200
rect 10945 -260 10965 -200
rect 11020 -260 11045 -200
rect 10870 -279 11045 -260
rect 10920 -280 11045 -279
rect 8120 -435 8425 -400
rect 9485 -360 9605 -340
rect 9485 -420 9525 -360
rect 9575 -420 9605 -360
rect 9485 -440 9605 -420
rect 7525 -450 7900 -445
rect 7525 -455 7565 -450
rect 9890 -500 9940 -290
rect 6845 -555 7475 -520
rect 9860 -510 9970 -500
rect 9860 -580 9870 -510
rect 9960 -580 9970 -510
rect 9860 -590 9970 -580
rect 10290 -610 10340 -280
rect 4840 -6750 10980 -610
<< viali >>
rect 4980 995 5000 1015
rect 4980 420 5005 440
rect 4925 360 4945 380
rect 5725 995 5745 1015
rect 6330 995 6350 1015
rect 5725 420 5750 440
rect 5675 360 5695 380
rect 7000 1770 7020 1790
rect 7000 1195 7025 1215
rect 6945 1135 6965 1155
rect 6995 1000 7015 1020
rect 7595 1770 7615 1790
rect 8635 1865 8660 1900
rect 8720 1865 8745 1900
rect 8905 1865 8930 1900
rect 8950 1865 8975 1900
rect 7595 1195 7620 1215
rect 7540 1135 7560 1155
rect 6330 420 6355 440
rect 6275 360 6295 380
rect 6995 425 7020 445
rect 6940 365 6960 385
rect 7590 1000 7610 1020
rect 7590 425 7615 445
rect 7535 365 7555 385
rect 9500 1710 9540 1750
rect 9560 1710 9600 1750
rect 9620 1710 9660 1750
rect 9680 1710 9720 1750
rect 9740 1710 9780 1750
rect 9800 1710 9840 1750
rect 9860 1710 9900 1750
rect 9920 1710 9960 1750
rect 9980 1710 10020 1750
rect 10040 1710 10080 1750
rect 10100 1710 10140 1750
rect 10160 1710 10200 1750
rect 10220 1710 10260 1750
rect 10280 1710 10320 1750
rect 10340 1710 10380 1750
rect 10400 1710 10440 1750
rect 10460 1710 10500 1750
rect 10520 1710 10560 1750
rect 9500 1650 9540 1690
rect 9560 1650 9600 1690
rect 9620 1650 9660 1690
rect 9680 1650 9720 1690
rect 9740 1650 9780 1690
rect 9800 1650 9840 1690
rect 9860 1650 9900 1690
rect 9920 1650 9960 1690
rect 9980 1650 10020 1690
rect 10040 1650 10080 1690
rect 10100 1650 10140 1690
rect 10160 1650 10200 1690
rect 10220 1650 10260 1690
rect 10280 1650 10320 1690
rect 10340 1650 10380 1690
rect 10400 1650 10440 1690
rect 10460 1650 10500 1690
rect 10520 1650 10560 1690
rect 8905 1565 8930 1600
rect 8950 1565 8975 1600
rect 7590 190 7610 210
rect 7590 -385 7615 -365
rect 9040 130 9130 205
rect 9130 130 9135 205
rect 10130 730 10195 795
rect 7535 -445 7555 -425
rect 10890 -260 10945 -200
rect 9525 -420 9575 -360
rect 9870 -580 9960 -510
<< metal1 >>
rect 8605 2175 8770 2300
rect 8855 2175 9020 2300
rect 8615 1900 8760 2175
rect 8615 1865 8635 1900
rect 8660 1865 8720 1900
rect 8745 1865 8760 1900
rect 8615 1845 8760 1865
rect 8865 1900 9010 2175
rect 9495 2080 9660 2205
rect 8865 1865 8905 1900
rect 8930 1865 8950 1900
rect 8975 1865 9010 1900
rect 8865 1845 9010 1865
rect 9505 1805 9650 2080
rect 10200 1805 10680 1810
rect 4895 1790 10680 1805
rect 4895 1770 7000 1790
rect 7020 1770 7595 1790
rect 7615 1770 10680 1790
rect 4895 1750 10680 1770
rect 4895 1030 4940 1750
rect 5565 1030 5610 1750
rect 6140 1030 6185 1750
rect 6845 1035 6890 1750
rect 6990 1215 7165 1220
rect 6990 1195 7000 1215
rect 7025 1195 7165 1215
rect 6990 1185 7165 1195
rect 6935 1160 6975 1165
rect 6935 1130 6940 1160
rect 6970 1130 6975 1160
rect 6935 1125 6975 1130
rect 4895 1015 5090 1030
rect 4895 995 4980 1015
rect 5000 995 5090 1015
rect 4895 975 5090 995
rect 5565 1015 5835 1030
rect 5565 995 5725 1015
rect 5745 995 5835 1015
rect 5565 975 5835 995
rect 6140 1015 6440 1030
rect 6140 995 6330 1015
rect 6350 995 6440 1015
rect 6140 975 6440 995
rect 6845 1020 7105 1035
rect 6845 1000 6995 1020
rect 7015 1000 7105 1020
rect 6845 975 7105 1000
rect 7130 450 7165 1185
rect 7440 1035 7485 1750
rect 9470 1710 9500 1750
rect 9540 1710 9560 1750
rect 9600 1710 9620 1750
rect 9660 1710 9680 1750
rect 9720 1710 9740 1750
rect 9780 1710 9800 1750
rect 9840 1710 9860 1750
rect 9900 1710 9920 1750
rect 9960 1710 9980 1750
rect 10020 1710 10040 1750
rect 10080 1710 10100 1750
rect 10140 1710 10160 1750
rect 10200 1710 10220 1750
rect 10260 1710 10280 1750
rect 10320 1710 10340 1750
rect 10380 1710 10400 1750
rect 10440 1710 10460 1750
rect 10500 1710 10520 1750
rect 10560 1710 10680 1750
rect 9470 1690 10680 1710
rect 9470 1650 9500 1690
rect 9540 1650 9560 1690
rect 9600 1650 9620 1690
rect 9660 1650 9680 1690
rect 9720 1650 9740 1690
rect 9780 1650 9800 1690
rect 9840 1650 9860 1690
rect 9900 1650 9920 1690
rect 9960 1650 9980 1690
rect 10020 1650 10040 1690
rect 10080 1650 10100 1690
rect 10140 1650 10160 1690
rect 10200 1650 10220 1690
rect 10260 1650 10280 1690
rect 10320 1650 10340 1690
rect 10380 1650 10400 1690
rect 10440 1650 10460 1690
rect 10500 1650 10520 1690
rect 10560 1650 10680 1690
rect 8895 1600 8985 1625
rect 9470 1620 10680 1650
rect 8895 1565 8905 1600
rect 8930 1565 8950 1600
rect 8975 1565 8985 1600
rect 7585 1215 7750 1220
rect 7585 1195 7595 1215
rect 7620 1195 7750 1215
rect 7585 1185 7750 1195
rect 7530 1160 7570 1165
rect 7530 1130 7535 1160
rect 7565 1130 7570 1160
rect 7530 1125 7570 1130
rect 7440 1030 7700 1035
rect 6985 445 7165 450
rect 4970 440 5140 445
rect 4970 420 4980 440
rect 5005 420 5140 440
rect 4970 410 5140 420
rect 5715 440 5885 445
rect 5715 420 5725 440
rect 5750 420 5885 440
rect 5715 410 5885 420
rect 6320 440 6490 445
rect 6320 420 6330 440
rect 6355 420 6490 440
rect 6320 410 6490 420
rect 6985 425 6995 445
rect 7020 425 7165 445
rect 6985 415 7165 425
rect 4915 385 4955 390
rect 4915 355 4920 385
rect 4950 355 4955 385
rect 4915 350 4955 355
rect 5105 -500 5140 410
rect 5665 385 5705 390
rect 5665 355 5670 385
rect 5700 355 5705 385
rect 5665 350 5705 355
rect 5850 -500 5885 410
rect 6265 385 6305 390
rect 6265 355 6270 385
rect 6300 355 6305 385
rect 6265 350 6305 355
rect 6455 -500 6490 410
rect 6930 390 6970 395
rect 6930 360 6935 390
rect 6965 360 6970 390
rect 6930 355 6970 360
rect 7130 -500 7165 415
rect 7435 1020 7700 1030
rect 7435 1000 7590 1020
rect 7610 1000 7700 1020
rect 7435 975 7700 1000
rect 7435 225 7480 975
rect 7715 450 7750 1185
rect 7580 445 7750 450
rect 7580 425 7590 445
rect 7615 425 7750 445
rect 7580 415 7750 425
rect 7525 390 7565 395
rect 7525 360 7530 390
rect 7560 360 7565 390
rect 7525 355 7565 360
rect 7435 210 7700 225
rect 7435 190 7590 210
rect 7610 190 7700 210
rect 7435 170 7700 190
rect 7715 -360 7750 415
rect 8895 220 8985 1565
rect 9890 795 10570 830
rect 9890 730 10130 795
rect 10195 730 10570 795
rect 9890 700 10570 730
rect 8895 205 9140 220
rect 8895 130 9040 205
rect 9135 130 9140 205
rect 8895 120 9140 130
rect 9890 -320 9980 700
rect 7580 -365 7750 -360
rect 7580 -385 7590 -365
rect 7615 -385 7750 -365
rect 7580 -395 7750 -385
rect 7525 -420 7565 -415
rect 7525 -450 7530 -420
rect 7560 -450 7565 -420
rect 7525 -455 7565 -450
rect 7715 -500 7750 -395
rect 9430 -360 9980 -320
rect 10505 -180 10570 700
rect 11205 -180 11300 -170
rect 10505 -200 11300 -180
rect 10505 -260 10890 -200
rect 10945 -260 11300 -200
rect 10505 -325 11300 -260
rect 11205 -335 11300 -325
rect 9430 -420 9525 -360
rect 9575 -410 9980 -360
rect 9575 -420 9650 -410
rect 9430 -500 9650 -420
rect 5105 -535 9650 -500
rect 9860 -510 9970 -500
rect 9860 -580 9870 -510
rect 9960 -580 9970 -510
rect 9860 -610 9970 -580
rect 4840 -6750 10980 -610
<< via1 >>
rect 6940 1155 6970 1160
rect 6940 1135 6945 1155
rect 6945 1135 6965 1155
rect 6965 1135 6970 1155
rect 6940 1130 6970 1135
rect 7535 1155 7565 1160
rect 7535 1135 7540 1155
rect 7540 1135 7560 1155
rect 7560 1135 7565 1155
rect 7535 1130 7565 1135
rect 4920 380 4950 385
rect 4920 360 4925 380
rect 4925 360 4945 380
rect 4945 360 4950 380
rect 4920 355 4950 360
rect 5670 380 5700 385
rect 5670 360 5675 380
rect 5675 360 5695 380
rect 5695 360 5700 380
rect 5670 355 5700 360
rect 6270 380 6300 385
rect 6270 360 6275 380
rect 6275 360 6295 380
rect 6295 360 6300 380
rect 6270 355 6300 360
rect 6935 385 6965 390
rect 6935 365 6940 385
rect 6940 365 6960 385
rect 6960 365 6965 385
rect 6935 360 6965 365
rect 7530 385 7560 390
rect 7530 365 7535 385
rect 7535 365 7555 385
rect 7555 365 7560 385
rect 7530 360 7560 365
rect 7530 -425 7560 -420
rect 7530 -445 7535 -425
rect 7535 -445 7555 -425
rect 7555 -445 7560 -425
rect 7530 -450 7560 -445
<< metal2 >>
rect 5900 2280 6000 2380
rect 6200 2280 6300 2380
rect 6500 2280 6600 2380
rect 6800 2280 6900 2380
rect 7100 2280 7200 2380
rect 7400 2280 7500 2380
rect 7700 2280 7800 2380
rect 8000 2280 8100 2380
rect 5930 2080 5970 2280
rect 5300 2035 5970 2080
rect 6230 2070 6270 2280
rect 5300 390 5340 2035
rect 6085 2025 6270 2070
rect 6540 2070 6580 2280
rect 6830 2070 6870 2280
rect 7130 2155 7175 2280
rect 7425 2255 7470 2280
rect 7425 2210 7595 2255
rect 7130 2110 7480 2155
rect 6540 2025 6780 2070
rect 6830 2025 7405 2070
rect 6085 390 6125 2025
rect 6740 390 6780 2025
rect 7365 1165 7405 2025
rect 7435 1915 7480 2110
rect 7550 2070 7595 2210
rect 7725 2155 7770 2280
rect 8025 2225 8070 2280
rect 8025 2190 8375 2225
rect 8025 2180 8380 2190
rect 7725 2110 8165 2155
rect 7550 2025 8045 2070
rect 6935 1160 7405 1165
rect 6935 1130 6940 1160
rect 6970 1130 7405 1160
rect 6935 1125 7405 1130
rect 7365 1120 7405 1125
rect 7440 395 7480 1915
rect 8005 1165 8045 2025
rect 7530 1160 8045 1165
rect 7530 1130 7535 1160
rect 7565 1130 8045 1160
rect 7530 1125 8045 1130
rect 8125 395 8165 2110
rect 4915 385 5340 390
rect 4915 355 4920 385
rect 4950 355 5340 385
rect 4915 350 5340 355
rect 5665 385 6125 390
rect 5665 355 5670 385
rect 5700 355 6125 385
rect 5665 350 6125 355
rect 6265 385 6780 390
rect 6265 355 6270 385
rect 6300 355 6780 385
rect 6930 390 7480 395
rect 6930 360 6935 390
rect 6965 360 7480 390
rect 6930 355 7480 360
rect 7525 390 8165 395
rect 7525 360 7530 390
rect 7560 360 8165 390
rect 7525 355 8165 360
rect 8335 2040 8380 2180
rect 6265 350 6780 355
rect 8335 -415 8375 2040
rect 7525 -420 8375 -415
rect 7525 -450 7530 -420
rect 7560 -450 8375 -420
rect 7525 -455 8375 -450
<< labels >>
flabel locali 9060 750 9170 850 0 FreeSans 800 0 0 0 A
flabel locali 9520 770 9570 820 0 FreeSans 800 0 0 0 B
flabel locali 9370 220 9420 250 0 FreeSans 800 0 0 0 C
flabel locali 9890 220 9940 270 0 FreeSans 800 0 0 0 D
flabel locali 10290 -440 10340 -390 0 FreeSans 800 0 0 0 E
flabel polycont 9040 260 9130 340 0 FreeSans 800 0 0 0 n0
flabel locali 8205 205 8240 395 0 FreeSans 800 0 0 0 n1
flabel locali 8205 910 8240 1050 0 FreeSans 800 0 0 0 n2
flabel locali 8205 1600 8240 1920 0 FreeSans 800 0 0 0 n3
flabel locali 7440 750 7475 980 0 FreeSans 800 0 0 0 n4
flabel locali 7440 -555 7475 -10 0 FreeSans 800 0 0 0 n5
flabel locali 6845 1600 6880 1920 0 FreeSans 800 0 0 0 n6
flabel locali 6140 -555 6175 0 0 FreeSans 800 0 0 0 n7
flabel locali 5440 1360 5565 1600 0 FreeSans 800 0 0 0 n8
flabel polycont 7860 220 7880 240 0 FreeSans 800 0 0 0 nc0
flabel polycont 7860 1030 7880 1050 0 FreeSans 800 0 0 0 nc1
flabel polycont 7865 1800 7885 1820 0 FreeSans 800 0 0 0 nc2
flabel polycont 7270 1800 7290 1820 0 FreeSans 800 0 0 0 nc3
flabel polycont 7265 1030 7285 1050 0 FreeSans 800 0 0 0 nc4
flabel polycont 6600 1025 6620 1045 0 FreeSans 800 0 0 0 nc5
flabel polycont 5995 1025 6015 1045 0 FreeSans 800 0 0 0 nc6
flabel polycont 5250 1025 5270 1045 0 FreeSans 800 0 0 0 nc7
flabel metal2 8000 2280 8100 2380 0 FreeSans 800 0 0 0 c0
flabel metal2 7700 2280 7800 2380 0 FreeSans 800 0 0 0 c1
flabel metal2 7400 2280 7500 2380 0 FreeSans 800 0 0 0 c2
flabel metal2 7100 2280 7200 2380 0 FreeSans 800 0 0 0 c4
flabel metal2 6800 2280 6900 2380 0 FreeSans 800 0 0 0 c3
flabel metal2 6500 2280 6600 2380 0 FreeSans 800 0 0 0 c5
flabel metal2 6200 2280 6300 2380 0 FreeSans 800 0 0 0 c6
flabel metal2 5900 2280 6000 2380 0 FreeSans 800 0 0 0 c7
flabel metal1 9495 2080 9660 2205 0 FreeSans 800 0 0 0 VD
flabel metal1 11205 -335 11300 -170 0 FreeSans 800 0 0 0 VS
flabel metal1 8605 2175 8770 2300 0 FreeSans 800 0 0 0 IN1
flabel metal1 8855 2175 9020 2300 0 FreeSans 800 0 0 0 IN2
flabel locali 11025 725 11130 825 0 FreeSans 800 0 0 0 OUT
<< end >>
