magic
tech sky130A
magscale 1 2
timestamp 1634602588
<< locali >>
rect 6745 2363 6779 2465
<< viali >>
rect 2513 18309 2547 18343
rect 11897 18241 11931 18275
rect 16129 18241 16163 18275
rect 2605 18037 2639 18071
rect 11713 18037 11747 18071
rect 15945 18037 15979 18071
rect 15853 17629 15887 17663
rect 15761 17493 15795 17527
rect 10885 5729 10919 5763
rect 9689 5661 9723 5695
rect 10609 5661 10643 5695
rect 10701 5661 10735 5695
rect 10977 5661 11011 5695
rect 12081 5661 12115 5695
rect 9505 5525 9539 5559
rect 10425 5525 10459 5559
rect 11897 5525 11931 5559
rect 9229 5321 9263 5355
rect 10701 5253 10735 5287
rect 12357 5185 12391 5219
rect 8493 5117 8527 5151
rect 8769 5117 8803 5151
rect 10977 5117 11011 5151
rect 12081 5117 12115 5151
rect 7021 4981 7055 5015
rect 6469 4641 6503 4675
rect 9597 4573 9631 4607
rect 12817 4573 12851 4607
rect 13093 4573 13127 4607
rect 14657 4573 14691 4607
rect 6745 4505 6779 4539
rect 8217 4437 8251 4471
rect 10885 4437 10919 4471
rect 14473 4437 14507 4471
rect 6837 4233 6871 4267
rect 7849 4233 7883 4267
rect 8493 4233 8527 4267
rect 7021 4097 7055 4131
rect 7113 4097 7147 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 9045 4097 9079 4131
rect 10333 4097 10367 4131
rect 10793 4097 10827 4131
rect 10885 4097 10919 4131
rect 11713 4097 11747 4131
rect 7297 4029 7331 4063
rect 10057 4029 10091 4063
rect 12541 4029 12575 4063
rect 12817 4029 12851 4063
rect 8953 3893 8987 3927
rect 11529 3893 11563 3927
rect 14289 3893 14323 3927
rect 12633 3689 12667 3723
rect 13093 3621 13127 3655
rect 10517 3553 10551 3587
rect 7021 3485 7055 3519
rect 7481 3485 7515 3519
rect 9597 3485 9631 3519
rect 10241 3485 10275 3519
rect 12817 3485 12851 3519
rect 12909 3485 12943 3519
rect 13185 3485 13219 3519
rect 8125 3417 8159 3451
rect 8309 3417 8343 3451
rect 14105 3417 14139 3451
rect 14289 3417 14323 3451
rect 5733 3349 5767 3383
rect 7665 3349 7699 3383
rect 9781 3349 9815 3383
rect 11989 3349 12023 3383
rect 8585 3145 8619 3179
rect 9321 3077 9355 3111
rect 9045 3009 9079 3043
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 11989 2941 12023 2975
rect 12265 2941 12299 2975
rect 10793 2805 10827 2839
rect 13737 2805 13771 2839
rect 6837 2601 6871 2635
rect 8401 2601 8435 2635
rect 10517 2601 10551 2635
rect 12265 2601 12299 2635
rect 14197 2601 14231 2635
rect 7297 2533 7331 2567
rect 14657 2533 14691 2567
rect 6745 2465 6779 2499
rect 7941 2465 7975 2499
rect 12725 2465 12759 2499
rect 1961 2397 1995 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 7113 2397 7147 2431
rect 7389 2397 7423 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 12449 2397 12483 2431
rect 12541 2397 12575 2431
rect 12817 2397 12851 2431
rect 14105 2397 14139 2431
rect 14381 2397 14415 2431
rect 14473 2397 14507 2431
rect 15945 2397 15979 2431
rect 1777 2329 1811 2363
rect 4169 2329 4203 2363
rect 5733 2329 5767 2363
rect 6745 2329 6779 2363
rect 9229 2329 9263 2363
rect 13277 2329 13311 2363
rect 13461 2329 13495 2363
rect 15117 2329 15151 2363
rect 15301 2329 15335 2363
rect 16129 2329 16163 2363
rect 5641 2261 5675 2295
<< metal1 >>
rect 1104 18522 17480 18544
rect 1104 18470 6408 18522
rect 6460 18470 6472 18522
rect 6524 18470 6536 18522
rect 6588 18470 6600 18522
rect 6652 18470 6664 18522
rect 6716 18470 11867 18522
rect 11919 18470 11931 18522
rect 11983 18470 11995 18522
rect 12047 18470 12059 18522
rect 12111 18470 12123 18522
rect 12175 18470 17480 18522
rect 1104 18448 17480 18470
rect 2314 18300 2320 18352
rect 2372 18340 2378 18352
rect 2501 18343 2559 18349
rect 2501 18340 2513 18343
rect 2372 18312 2513 18340
rect 2372 18300 2378 18312
rect 2501 18309 2513 18312
rect 2547 18309 2559 18343
rect 2501 18303 2559 18309
rect 11606 18232 11612 18284
rect 11664 18272 11670 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11664 18244 11897 18272
rect 11664 18232 11670 18244
rect 11885 18241 11897 18244
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16206 18272 16212 18284
rect 16163 18244 16212 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 2593 18071 2651 18077
rect 2593 18037 2605 18071
rect 2639 18068 2651 18071
rect 10594 18068 10600 18080
rect 2639 18040 10600 18068
rect 2639 18037 2651 18040
rect 2593 18031 2651 18037
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15896 18040 15945 18068
rect 15896 18028 15902 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 1104 17978 17480 18000
rect 1104 17926 3679 17978
rect 3731 17926 3743 17978
rect 3795 17926 3807 17978
rect 3859 17926 3871 17978
rect 3923 17926 3935 17978
rect 3987 17926 9138 17978
rect 9190 17926 9202 17978
rect 9254 17926 9266 17978
rect 9318 17926 9330 17978
rect 9382 17926 9394 17978
rect 9446 17926 14596 17978
rect 14648 17926 14660 17978
rect 14712 17926 14724 17978
rect 14776 17926 14788 17978
rect 14840 17926 14852 17978
rect 14904 17926 17480 17978
rect 1104 17904 17480 17926
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 9582 17864 9588 17876
rect 6972 17836 9588 17864
rect 6972 17824 6978 17836
rect 9582 17824 9588 17836
rect 9640 17824 9646 17876
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 15746 17524 15752 17536
rect 15707 17496 15752 17524
rect 15746 17484 15752 17496
rect 15804 17484 15810 17536
rect 1104 17434 17480 17456
rect 1104 17382 6408 17434
rect 6460 17382 6472 17434
rect 6524 17382 6536 17434
rect 6588 17382 6600 17434
rect 6652 17382 6664 17434
rect 6716 17382 11867 17434
rect 11919 17382 11931 17434
rect 11983 17382 11995 17434
rect 12047 17382 12059 17434
rect 12111 17382 12123 17434
rect 12175 17382 17480 17434
rect 1104 17360 17480 17382
rect 1104 16890 17480 16912
rect 1104 16838 3679 16890
rect 3731 16838 3743 16890
rect 3795 16838 3807 16890
rect 3859 16838 3871 16890
rect 3923 16838 3935 16890
rect 3987 16838 9138 16890
rect 9190 16838 9202 16890
rect 9254 16838 9266 16890
rect 9318 16838 9330 16890
rect 9382 16838 9394 16890
rect 9446 16838 14596 16890
rect 14648 16838 14660 16890
rect 14712 16838 14724 16890
rect 14776 16838 14788 16890
rect 14840 16838 14852 16890
rect 14904 16838 17480 16890
rect 1104 16816 17480 16838
rect 1104 16346 17480 16368
rect 1104 16294 6408 16346
rect 6460 16294 6472 16346
rect 6524 16294 6536 16346
rect 6588 16294 6600 16346
rect 6652 16294 6664 16346
rect 6716 16294 11867 16346
rect 11919 16294 11931 16346
rect 11983 16294 11995 16346
rect 12047 16294 12059 16346
rect 12111 16294 12123 16346
rect 12175 16294 17480 16346
rect 1104 16272 17480 16294
rect 1104 15802 17480 15824
rect 1104 15750 3679 15802
rect 3731 15750 3743 15802
rect 3795 15750 3807 15802
rect 3859 15750 3871 15802
rect 3923 15750 3935 15802
rect 3987 15750 9138 15802
rect 9190 15750 9202 15802
rect 9254 15750 9266 15802
rect 9318 15750 9330 15802
rect 9382 15750 9394 15802
rect 9446 15750 14596 15802
rect 14648 15750 14660 15802
rect 14712 15750 14724 15802
rect 14776 15750 14788 15802
rect 14840 15750 14852 15802
rect 14904 15750 17480 15802
rect 1104 15728 17480 15750
rect 1104 15258 17480 15280
rect 1104 15206 6408 15258
rect 6460 15206 6472 15258
rect 6524 15206 6536 15258
rect 6588 15206 6600 15258
rect 6652 15206 6664 15258
rect 6716 15206 11867 15258
rect 11919 15206 11931 15258
rect 11983 15206 11995 15258
rect 12047 15206 12059 15258
rect 12111 15206 12123 15258
rect 12175 15206 17480 15258
rect 1104 15184 17480 15206
rect 1104 14714 17480 14736
rect 1104 14662 3679 14714
rect 3731 14662 3743 14714
rect 3795 14662 3807 14714
rect 3859 14662 3871 14714
rect 3923 14662 3935 14714
rect 3987 14662 9138 14714
rect 9190 14662 9202 14714
rect 9254 14662 9266 14714
rect 9318 14662 9330 14714
rect 9382 14662 9394 14714
rect 9446 14662 14596 14714
rect 14648 14662 14660 14714
rect 14712 14662 14724 14714
rect 14776 14662 14788 14714
rect 14840 14662 14852 14714
rect 14904 14662 17480 14714
rect 1104 14640 17480 14662
rect 1104 14170 17480 14192
rect 1104 14118 6408 14170
rect 6460 14118 6472 14170
rect 6524 14118 6536 14170
rect 6588 14118 6600 14170
rect 6652 14118 6664 14170
rect 6716 14118 11867 14170
rect 11919 14118 11931 14170
rect 11983 14118 11995 14170
rect 12047 14118 12059 14170
rect 12111 14118 12123 14170
rect 12175 14118 17480 14170
rect 1104 14096 17480 14118
rect 1104 13626 17480 13648
rect 1104 13574 3679 13626
rect 3731 13574 3743 13626
rect 3795 13574 3807 13626
rect 3859 13574 3871 13626
rect 3923 13574 3935 13626
rect 3987 13574 9138 13626
rect 9190 13574 9202 13626
rect 9254 13574 9266 13626
rect 9318 13574 9330 13626
rect 9382 13574 9394 13626
rect 9446 13574 14596 13626
rect 14648 13574 14660 13626
rect 14712 13574 14724 13626
rect 14776 13574 14788 13626
rect 14840 13574 14852 13626
rect 14904 13574 17480 13626
rect 1104 13552 17480 13574
rect 1104 13082 17480 13104
rect 1104 13030 6408 13082
rect 6460 13030 6472 13082
rect 6524 13030 6536 13082
rect 6588 13030 6600 13082
rect 6652 13030 6664 13082
rect 6716 13030 11867 13082
rect 11919 13030 11931 13082
rect 11983 13030 11995 13082
rect 12047 13030 12059 13082
rect 12111 13030 12123 13082
rect 12175 13030 17480 13082
rect 1104 13008 17480 13030
rect 1104 12538 17480 12560
rect 1104 12486 3679 12538
rect 3731 12486 3743 12538
rect 3795 12486 3807 12538
rect 3859 12486 3871 12538
rect 3923 12486 3935 12538
rect 3987 12486 9138 12538
rect 9190 12486 9202 12538
rect 9254 12486 9266 12538
rect 9318 12486 9330 12538
rect 9382 12486 9394 12538
rect 9446 12486 14596 12538
rect 14648 12486 14660 12538
rect 14712 12486 14724 12538
rect 14776 12486 14788 12538
rect 14840 12486 14852 12538
rect 14904 12486 17480 12538
rect 1104 12464 17480 12486
rect 1104 11994 17480 12016
rect 1104 11942 6408 11994
rect 6460 11942 6472 11994
rect 6524 11942 6536 11994
rect 6588 11942 6600 11994
rect 6652 11942 6664 11994
rect 6716 11942 11867 11994
rect 11919 11942 11931 11994
rect 11983 11942 11995 11994
rect 12047 11942 12059 11994
rect 12111 11942 12123 11994
rect 12175 11942 17480 11994
rect 1104 11920 17480 11942
rect 1104 11450 17480 11472
rect 1104 11398 3679 11450
rect 3731 11398 3743 11450
rect 3795 11398 3807 11450
rect 3859 11398 3871 11450
rect 3923 11398 3935 11450
rect 3987 11398 9138 11450
rect 9190 11398 9202 11450
rect 9254 11398 9266 11450
rect 9318 11398 9330 11450
rect 9382 11398 9394 11450
rect 9446 11398 14596 11450
rect 14648 11398 14660 11450
rect 14712 11398 14724 11450
rect 14776 11398 14788 11450
rect 14840 11398 14852 11450
rect 14904 11398 17480 11450
rect 1104 11376 17480 11398
rect 1104 10906 17480 10928
rect 1104 10854 6408 10906
rect 6460 10854 6472 10906
rect 6524 10854 6536 10906
rect 6588 10854 6600 10906
rect 6652 10854 6664 10906
rect 6716 10854 11867 10906
rect 11919 10854 11931 10906
rect 11983 10854 11995 10906
rect 12047 10854 12059 10906
rect 12111 10854 12123 10906
rect 12175 10854 17480 10906
rect 1104 10832 17480 10854
rect 1104 10362 17480 10384
rect 1104 10310 3679 10362
rect 3731 10310 3743 10362
rect 3795 10310 3807 10362
rect 3859 10310 3871 10362
rect 3923 10310 3935 10362
rect 3987 10310 9138 10362
rect 9190 10310 9202 10362
rect 9254 10310 9266 10362
rect 9318 10310 9330 10362
rect 9382 10310 9394 10362
rect 9446 10310 14596 10362
rect 14648 10310 14660 10362
rect 14712 10310 14724 10362
rect 14776 10310 14788 10362
rect 14840 10310 14852 10362
rect 14904 10310 17480 10362
rect 1104 10288 17480 10310
rect 1104 9818 17480 9840
rect 1104 9766 6408 9818
rect 6460 9766 6472 9818
rect 6524 9766 6536 9818
rect 6588 9766 6600 9818
rect 6652 9766 6664 9818
rect 6716 9766 11867 9818
rect 11919 9766 11931 9818
rect 11983 9766 11995 9818
rect 12047 9766 12059 9818
rect 12111 9766 12123 9818
rect 12175 9766 17480 9818
rect 1104 9744 17480 9766
rect 1104 9274 17480 9296
rect 1104 9222 3679 9274
rect 3731 9222 3743 9274
rect 3795 9222 3807 9274
rect 3859 9222 3871 9274
rect 3923 9222 3935 9274
rect 3987 9222 9138 9274
rect 9190 9222 9202 9274
rect 9254 9222 9266 9274
rect 9318 9222 9330 9274
rect 9382 9222 9394 9274
rect 9446 9222 14596 9274
rect 14648 9222 14660 9274
rect 14712 9222 14724 9274
rect 14776 9222 14788 9274
rect 14840 9222 14852 9274
rect 14904 9222 17480 9274
rect 1104 9200 17480 9222
rect 1104 8730 17480 8752
rect 1104 8678 6408 8730
rect 6460 8678 6472 8730
rect 6524 8678 6536 8730
rect 6588 8678 6600 8730
rect 6652 8678 6664 8730
rect 6716 8678 11867 8730
rect 11919 8678 11931 8730
rect 11983 8678 11995 8730
rect 12047 8678 12059 8730
rect 12111 8678 12123 8730
rect 12175 8678 17480 8730
rect 1104 8656 17480 8678
rect 1104 8186 17480 8208
rect 1104 8134 3679 8186
rect 3731 8134 3743 8186
rect 3795 8134 3807 8186
rect 3859 8134 3871 8186
rect 3923 8134 3935 8186
rect 3987 8134 9138 8186
rect 9190 8134 9202 8186
rect 9254 8134 9266 8186
rect 9318 8134 9330 8186
rect 9382 8134 9394 8186
rect 9446 8134 14596 8186
rect 14648 8134 14660 8186
rect 14712 8134 14724 8186
rect 14776 8134 14788 8186
rect 14840 8134 14852 8186
rect 14904 8134 17480 8186
rect 1104 8112 17480 8134
rect 1104 7642 17480 7664
rect 1104 7590 6408 7642
rect 6460 7590 6472 7642
rect 6524 7590 6536 7642
rect 6588 7590 6600 7642
rect 6652 7590 6664 7642
rect 6716 7590 11867 7642
rect 11919 7590 11931 7642
rect 11983 7590 11995 7642
rect 12047 7590 12059 7642
rect 12111 7590 12123 7642
rect 12175 7590 17480 7642
rect 1104 7568 17480 7590
rect 1104 7098 17480 7120
rect 1104 7046 3679 7098
rect 3731 7046 3743 7098
rect 3795 7046 3807 7098
rect 3859 7046 3871 7098
rect 3923 7046 3935 7098
rect 3987 7046 9138 7098
rect 9190 7046 9202 7098
rect 9254 7046 9266 7098
rect 9318 7046 9330 7098
rect 9382 7046 9394 7098
rect 9446 7046 14596 7098
rect 14648 7046 14660 7098
rect 14712 7046 14724 7098
rect 14776 7046 14788 7098
rect 14840 7046 14852 7098
rect 14904 7046 17480 7098
rect 1104 7024 17480 7046
rect 1104 6554 17480 6576
rect 1104 6502 6408 6554
rect 6460 6502 6472 6554
rect 6524 6502 6536 6554
rect 6588 6502 6600 6554
rect 6652 6502 6664 6554
rect 6716 6502 11867 6554
rect 11919 6502 11931 6554
rect 11983 6502 11995 6554
rect 12047 6502 12059 6554
rect 12111 6502 12123 6554
rect 12175 6502 17480 6554
rect 1104 6480 17480 6502
rect 1104 6010 17480 6032
rect 1104 5958 3679 6010
rect 3731 5958 3743 6010
rect 3795 5958 3807 6010
rect 3859 5958 3871 6010
rect 3923 5958 3935 6010
rect 3987 5958 9138 6010
rect 9190 5958 9202 6010
rect 9254 5958 9266 6010
rect 9318 5958 9330 6010
rect 9382 5958 9394 6010
rect 9446 5958 14596 6010
rect 14648 5958 14660 6010
rect 14712 5958 14724 6010
rect 14776 5958 14788 6010
rect 14840 5958 14852 6010
rect 14904 5958 17480 6010
rect 1104 5936 17480 5958
rect 9692 5800 11468 5828
rect 9692 5701 9720 5800
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 9824 5732 10885 5760
rect 9824 5720 9830 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10873 5723 10931 5729
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 10594 5692 10600 5704
rect 10555 5664 10600 5692
rect 9677 5655 9735 5661
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11054 5692 11060 5704
rect 11011 5664 11060 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 10704 5624 10732 5655
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11440 5692 11468 5800
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11440 5664 12081 5692
rect 12069 5661 12081 5664
rect 12115 5692 12127 5695
rect 13078 5692 13084 5704
rect 12115 5664 13084 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 11698 5624 11704 5636
rect 10704 5596 11704 5624
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9456 5528 9505 5556
rect 9456 5516 9462 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 10410 5556 10416 5568
rect 10371 5528 10416 5556
rect 9493 5519 9551 5525
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11790 5516 11796 5568
rect 11848 5556 11854 5568
rect 11885 5559 11943 5565
rect 11885 5556 11897 5559
rect 11848 5528 11897 5556
rect 11848 5516 11854 5528
rect 11885 5525 11897 5528
rect 11931 5525 11943 5559
rect 11885 5519 11943 5525
rect 1104 5466 17480 5488
rect 1104 5414 6408 5466
rect 6460 5414 6472 5466
rect 6524 5414 6536 5466
rect 6588 5414 6600 5466
rect 6652 5414 6664 5466
rect 6716 5414 11867 5466
rect 11919 5414 11931 5466
rect 11983 5414 11995 5466
rect 12047 5414 12059 5466
rect 12111 5414 12123 5466
rect 12175 5414 17480 5466
rect 1104 5392 17480 5414
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 9217 5355 9275 5361
rect 9217 5352 9229 5355
rect 8904 5324 9229 5352
rect 8904 5312 8910 5324
rect 9217 5321 9229 5324
rect 9263 5352 9275 5355
rect 9766 5352 9772 5364
rect 9263 5324 9772 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 11790 5352 11796 5364
rect 10244 5324 11796 5352
rect 9398 5284 9404 5296
rect 8050 5256 9404 5284
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 10244 5270 10272 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 10410 5244 10416 5296
rect 10468 5284 10474 5296
rect 10689 5287 10747 5293
rect 10689 5284 10701 5287
rect 10468 5256 10701 5284
rect 10468 5244 10474 5256
rect 10689 5253 10701 5256
rect 10735 5253 10747 5287
rect 10689 5247 10747 5253
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 11112 5188 12357 5216
rect 11112 5176 11118 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 8478 5148 8484 5160
rect 8439 5120 8484 5148
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 8754 5148 8760 5160
rect 8715 5120 8760 5148
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 10962 5148 10968 5160
rect 10923 5120 10968 5148
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11790 5108 11796 5160
rect 11848 5148 11854 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11848 5120 12081 5148
rect 11848 5108 11854 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7009 5015 7067 5021
rect 7009 5012 7021 5015
rect 6972 4984 7021 5012
rect 6972 4972 6978 4984
rect 7009 4981 7021 4984
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 1104 4922 17480 4944
rect 1104 4870 3679 4922
rect 3731 4870 3743 4922
rect 3795 4870 3807 4922
rect 3859 4870 3871 4922
rect 3923 4870 3935 4922
rect 3987 4870 9138 4922
rect 9190 4870 9202 4922
rect 9254 4870 9266 4922
rect 9318 4870 9330 4922
rect 9382 4870 9394 4922
rect 9446 4870 14596 4922
rect 14648 4870 14660 4922
rect 14712 4870 14724 4922
rect 14776 4870 14788 4922
rect 14840 4870 14852 4922
rect 14904 4870 17480 4922
rect 1104 4848 17480 4870
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 8754 4672 8760 4684
rect 6503 4644 8760 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 7834 4564 7840 4616
rect 7892 4564 7898 4616
rect 9582 4604 9588 4616
rect 9543 4576 9588 4604
rect 9582 4564 9588 4576
rect 9640 4564 9646 4616
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 12894 4604 12900 4616
rect 12851 4576 12900 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13078 4604 13084 4616
rect 12991 4576 13084 4604
rect 13078 4564 13084 4576
rect 13136 4604 13142 4616
rect 14645 4607 14703 4613
rect 14645 4604 14657 4607
rect 13136 4576 14657 4604
rect 13136 4564 13142 4576
rect 14645 4573 14657 4576
rect 14691 4604 14703 4607
rect 15746 4604 15752 4616
rect 14691 4576 15752 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 6730 4536 6736 4548
rect 6691 4508 6736 4536
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 9732 4440 10885 4468
rect 9732 4428 9738 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 14458 4468 14464 4480
rect 14419 4440 14464 4468
rect 10873 4431 10931 4437
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 1104 4378 17480 4400
rect 1104 4326 6408 4378
rect 6460 4326 6472 4378
rect 6524 4326 6536 4378
rect 6588 4326 6600 4378
rect 6652 4326 6664 4378
rect 6716 4326 11867 4378
rect 11919 4326 11931 4378
rect 11983 4326 11995 4378
rect 12047 4326 12059 4378
rect 12111 4326 12123 4378
rect 12175 4326 17480 4378
rect 1104 4304 17480 4326
rect 6730 4224 6736 4276
rect 6788 4264 6794 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6788 4236 6837 4264
rect 6788 4224 6794 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 7834 4264 7840 4276
rect 7795 4236 7840 4264
rect 6825 4227 6883 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8478 4264 8484 4276
rect 8439 4236 8484 4264
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 6914 4156 6920 4208
rect 6972 4196 6978 4208
rect 6972 4168 7144 4196
rect 6972 4156 6978 4168
rect 7116 4137 7144 4168
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 12894 4196 12900 4208
rect 8352 4168 8800 4196
rect 8352 4156 8358 4168
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4097 7159 4131
rect 7101 4091 7159 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7834 4128 7840 4140
rect 7423 4100 7840 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7024 3992 7052 4091
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 8018 4128 8024 4140
rect 7979 4100 8024 4128
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8772 4137 8800 4168
rect 8956 4168 9168 4196
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4128 8815 4131
rect 8846 4128 8852 4140
rect 8803 4100 8852 4128
rect 8803 4097 8815 4100
rect 8757 4091 8815 4097
rect 7282 4060 7288 4072
rect 7195 4032 7288 4060
rect 7282 4020 7288 4032
rect 7340 4060 7346 4072
rect 8202 4060 8208 4072
rect 7340 4032 8208 4060
rect 7340 4020 7346 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8680 4060 8708 4091
rect 8846 4088 8852 4100
rect 8904 4088 8910 4140
rect 8956 4060 8984 4168
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4097 9091 4131
rect 9140 4128 9168 4168
rect 12452 4168 12900 4196
rect 10321 4131 10379 4137
rect 10321 4128 10333 4131
rect 9140 4100 10333 4128
rect 9033 4091 9091 4097
rect 10321 4097 10333 4100
rect 10367 4128 10379 4131
rect 10594 4128 10600 4140
rect 10367 4100 10600 4128
rect 10367 4097 10379 4100
rect 10321 4091 10379 4097
rect 8680 4032 8984 4060
rect 8680 3992 8708 4032
rect 9048 4004 9076 4091
rect 10594 4088 10600 4100
rect 10652 4128 10658 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10652 4100 10793 4128
rect 10652 4088 10658 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 11054 4128 11060 4140
rect 10919 4100 11060 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12452 4128 12480 4168
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 14458 4196 14464 4208
rect 14030 4168 14464 4196
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 11747 4100 12480 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 10042 4060 10048 4072
rect 10003 4032 10048 4060
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 11790 4060 11796 4072
rect 10152 4032 11796 4060
rect 9030 3992 9036 4004
rect 7024 3964 8708 3992
rect 8943 3964 9036 3992
rect 9030 3952 9036 3964
rect 9088 3992 9094 4004
rect 10152 3992 10180 4032
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4029 12587 4063
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12529 4023 12587 4029
rect 9088 3964 10180 3992
rect 9088 3952 9094 3964
rect 10226 3952 10232 4004
rect 10284 3992 10290 4004
rect 10962 3992 10968 4004
rect 10284 3964 10968 3992
rect 10284 3952 10290 3964
rect 10962 3952 10968 3964
rect 11020 3992 11026 4004
rect 12544 3992 12572 4023
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 11020 3964 12572 3992
rect 11020 3952 11026 3964
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 6972 3896 8953 3924
rect 6972 3884 6978 3896
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 8941 3887 8999 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 14277 3927 14335 3933
rect 14277 3893 14289 3927
rect 14323 3924 14335 3927
rect 14918 3924 14924 3936
rect 14323 3896 14924 3924
rect 14323 3893 14335 3896
rect 14277 3887 14335 3893
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 1104 3834 17480 3856
rect 1104 3782 3679 3834
rect 3731 3782 3743 3834
rect 3795 3782 3807 3834
rect 3859 3782 3871 3834
rect 3923 3782 3935 3834
rect 3987 3782 9138 3834
rect 9190 3782 9202 3834
rect 9254 3782 9266 3834
rect 9318 3782 9330 3834
rect 9382 3782 9394 3834
rect 9446 3782 14596 3834
rect 14648 3782 14660 3834
rect 14712 3782 14724 3834
rect 14776 3782 14788 3834
rect 14840 3782 14852 3834
rect 14904 3782 17480 3834
rect 1104 3760 17480 3782
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 9030 3720 9036 3732
rect 7892 3692 9036 3720
rect 7892 3680 7898 3692
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 12250 3720 12256 3732
rect 11112 3692 12256 3720
rect 11112 3680 11118 3692
rect 12250 3680 12256 3692
rect 12308 3720 12314 3732
rect 12621 3723 12679 3729
rect 12308 3692 12434 3720
rect 12308 3680 12314 3692
rect 9674 3652 9680 3664
rect 7024 3624 9680 3652
rect 7024 3525 7052 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 12406 3652 12434 3692
rect 12621 3689 12633 3723
rect 12667 3720 12679 3723
rect 12802 3720 12808 3732
rect 12667 3692 12808 3720
rect 12667 3689 12679 3692
rect 12621 3683 12679 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 13081 3655 13139 3661
rect 13081 3652 13093 3655
rect 12406 3624 13093 3652
rect 13081 3621 13093 3624
rect 13127 3621 13139 3655
rect 13081 3615 13139 3621
rect 8018 3544 8024 3596
rect 8076 3544 8082 3596
rect 10505 3587 10563 3593
rect 10505 3553 10517 3587
rect 10551 3584 10563 3587
rect 12342 3584 12348 3596
rect 10551 3556 12348 3584
rect 10551 3553 10563 3556
rect 10505 3547 10563 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12492 3556 12940 3584
rect 12492 3544 12498 3556
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3516 7527 3519
rect 8036 3516 8064 3544
rect 9585 3519 9643 3525
rect 9585 3516 9597 3519
rect 7515 3488 9597 3516
rect 7515 3485 7527 3488
rect 7469 3479 7527 3485
rect 9585 3485 9597 3488
rect 9631 3516 9643 3519
rect 10226 3516 10232 3528
rect 9631 3488 9904 3516
rect 10187 3488 10232 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 8076 3420 8125 3448
rect 8076 3408 8082 3420
rect 8113 3417 8125 3420
rect 8159 3417 8171 3451
rect 8113 3411 8171 3417
rect 8297 3451 8355 3457
rect 8297 3417 8309 3451
rect 8343 3448 8355 3451
rect 8570 3448 8576 3460
rect 8343 3420 8576 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 8570 3408 8576 3420
rect 8628 3408 8634 3460
rect 5718 3380 5724 3392
rect 5679 3352 5724 3380
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 7650 3380 7656 3392
rect 7611 3352 7656 3380
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 9766 3380 9772 3392
rect 9727 3352 9772 3380
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 9876 3380 9904 3488
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 12802 3516 12808 3528
rect 12763 3488 12808 3516
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 12912 3525 12940 3556
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13078 3516 13084 3528
rect 12943 3488 13084 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 14918 3516 14924 3528
rect 13219 3488 14924 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 11514 3408 11520 3460
rect 11572 3408 11578 3460
rect 11808 3420 12664 3448
rect 11808 3380 11836 3420
rect 9876 3352 11836 3380
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3380 12035 3383
rect 12526 3380 12532 3392
rect 12023 3352 12532 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12636 3380 12664 3420
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 12768 3420 14105 3448
rect 12768 3408 12774 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14274 3448 14280 3460
rect 14235 3420 14280 3448
rect 14093 3411 14151 3417
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 12894 3380 12900 3392
rect 12636 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 1104 3290 17480 3312
rect 1104 3238 6408 3290
rect 6460 3238 6472 3290
rect 6524 3238 6536 3290
rect 6588 3238 6600 3290
rect 6652 3238 6664 3290
rect 6716 3238 11867 3290
rect 11919 3238 11931 3290
rect 11983 3238 11995 3290
rect 12047 3238 12059 3290
rect 12111 3238 12123 3290
rect 12175 3238 17480 3290
rect 1104 3216 17480 3238
rect 8570 3176 8576 3188
rect 8531 3148 8576 3176
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 7650 3068 7656 3120
rect 7708 3068 7714 3120
rect 8386 3068 8392 3120
rect 8444 3108 8450 3120
rect 9309 3111 9367 3117
rect 9309 3108 9321 3111
rect 8444 3080 9321 3108
rect 8444 3068 8450 3080
rect 9309 3077 9321 3080
rect 9355 3077 9367 3111
rect 9309 3071 9367 3077
rect 9766 3068 9772 3120
rect 9824 3068 9830 3120
rect 12894 3068 12900 3120
rect 12952 3068 12958 3120
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8812 3012 9045 3040
rect 8812 3000 8818 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 5718 2932 5724 2984
rect 5776 2972 5782 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5776 2944 6837 2972
rect 5776 2932 5782 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 6825 2935 6883 2941
rect 6840 2836 6868 2935
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 10318 2932 10324 2984
rect 10376 2972 10382 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 10376 2944 11989 2972
rect 10376 2932 10382 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 12250 2972 12256 2984
rect 12211 2944 12256 2972
rect 11977 2935 12035 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 8754 2836 8760 2848
rect 6840 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 10778 2836 10784 2848
rect 10739 2808 10784 2836
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 13722 2836 13728 2848
rect 13683 2808 13728 2836
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 1104 2746 17480 2768
rect 1104 2694 3679 2746
rect 3731 2694 3743 2746
rect 3795 2694 3807 2746
rect 3859 2694 3871 2746
rect 3923 2694 3935 2746
rect 3987 2694 9138 2746
rect 9190 2694 9202 2746
rect 9254 2694 9266 2746
rect 9318 2694 9330 2746
rect 9382 2694 9394 2746
rect 9446 2694 14596 2746
rect 14648 2694 14660 2746
rect 14712 2694 14724 2746
rect 14776 2694 14788 2746
rect 14840 2694 14852 2746
rect 14904 2694 17480 2746
rect 1104 2672 17480 2694
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7098 2632 7104 2644
rect 6871 2604 7104 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 8202 2632 8208 2644
rect 7208 2604 8208 2632
rect 7208 2564 7236 2604
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10505 2635 10563 2641
rect 10505 2632 10517 2635
rect 10284 2604 10517 2632
rect 10284 2592 10290 2604
rect 10505 2601 10517 2604
rect 10551 2601 10563 2635
rect 12250 2632 12256 2644
rect 12211 2604 12256 2632
rect 10505 2595 10563 2601
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12526 2592 12532 2644
rect 12584 2632 12590 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 12584 2604 14197 2632
rect 12584 2592 12590 2604
rect 14185 2601 14197 2604
rect 14231 2632 14243 2635
rect 14274 2632 14280 2644
rect 14231 2604 14280 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 1964 2536 7236 2564
rect 7285 2567 7343 2573
rect 1964 2437 1992 2536
rect 7285 2533 7297 2567
rect 7331 2564 7343 2567
rect 8570 2564 8576 2576
rect 7331 2536 8576 2564
rect 7331 2533 7343 2536
rect 7285 2527 7343 2533
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7929 2499 7987 2505
rect 6779 2468 7144 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 6914 2428 6920 2440
rect 4387 2400 6920 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7116 2437 7144 2468
rect 7929 2465 7941 2499
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2428 7159 2431
rect 7282 2428 7288 2440
rect 7147 2400 7288 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 1118 2320 1124 2372
rect 1176 2360 1182 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1176 2332 1777 2360
rect 1176 2320 1182 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 3418 2320 3424 2372
rect 3476 2360 3482 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 3476 2332 4169 2360
rect 3476 2320 3482 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 5721 2363 5779 2369
rect 5721 2329 5733 2363
rect 5767 2360 5779 2363
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 5767 2332 6745 2360
rect 5767 2329 5779 2332
rect 5721 2323 5779 2329
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 6733 2323 6791 2329
rect 5626 2292 5632 2304
rect 5587 2264 5632 2292
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 7024 2292 7052 2391
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2428 7435 2431
rect 7834 2428 7840 2440
rect 7423 2400 7840 2428
rect 7423 2397 7435 2400
rect 7377 2391 7435 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7944 2360 7972 2459
rect 8036 2428 8064 2536
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 14645 2567 14703 2573
rect 14645 2564 14657 2567
rect 12400 2536 14657 2564
rect 12400 2524 12406 2536
rect 14645 2533 14657 2536
rect 14691 2533 14703 2567
rect 14645 2527 14703 2533
rect 10042 2496 10048 2508
rect 8220 2468 10048 2496
rect 8220 2440 8248 2468
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 10100 2468 10916 2496
rect 10100 2456 10106 2468
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 8036 2400 8125 2428
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 10778 2428 10784 2440
rect 8260 2400 8305 2428
rect 9140 2400 10784 2428
rect 8260 2388 8266 2400
rect 9140 2360 9168 2400
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 10888 2428 10916 2468
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12216 2468 12725 2496
rect 12216 2456 12222 2468
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 13078 2456 13084 2508
rect 13136 2496 13142 2508
rect 13136 2468 14504 2496
rect 13136 2456 13142 2468
rect 12434 2428 12440 2440
rect 10888 2400 12440 2428
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12584 2400 12629 2428
rect 12584 2388 12590 2400
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 13354 2428 13360 2440
rect 12860 2400 13360 2428
rect 12860 2388 12866 2400
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14476 2437 14504 2468
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 7944 2332 9168 2360
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2360 9275 2363
rect 9674 2360 9680 2372
rect 9263 2332 9680 2360
rect 9263 2329 9275 2332
rect 9217 2323 9275 2329
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 10468 2332 13277 2360
rect 10468 2320 10474 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 13449 2363 13507 2369
rect 13449 2329 13461 2363
rect 13495 2360 13507 2363
rect 14384 2360 14412 2391
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 14976 2400 15945 2428
rect 14976 2388 14982 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 13495 2332 14412 2360
rect 13495 2329 13507 2332
rect 13449 2323 13507 2329
rect 8202 2292 8208 2304
rect 7024 2264 8208 2292
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 10778 2252 10784 2304
rect 10836 2292 10842 2304
rect 13464 2292 13492 2323
rect 15010 2320 15016 2372
rect 15068 2360 15074 2372
rect 15105 2363 15163 2369
rect 15105 2360 15117 2363
rect 15068 2332 15117 2360
rect 15068 2320 15074 2332
rect 15105 2329 15117 2332
rect 15151 2329 15163 2363
rect 15105 2323 15163 2329
rect 15289 2363 15347 2369
rect 15289 2329 15301 2363
rect 15335 2329 15347 2363
rect 15289 2323 15347 2329
rect 16117 2363 16175 2369
rect 16117 2329 16129 2363
rect 16163 2360 16175 2363
rect 17310 2360 17316 2372
rect 16163 2332 17316 2360
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 10836 2264 13492 2292
rect 10836 2252 10842 2264
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 15304 2292 15332 2323
rect 17310 2320 17316 2332
rect 17368 2320 17374 2372
rect 13780 2264 15332 2292
rect 13780 2252 13786 2264
rect 1104 2202 17480 2224
rect 1104 2150 6408 2202
rect 6460 2150 6472 2202
rect 6524 2150 6536 2202
rect 6588 2150 6600 2202
rect 6652 2150 6664 2202
rect 6716 2150 11867 2202
rect 11919 2150 11931 2202
rect 11983 2150 11995 2202
rect 12047 2150 12059 2202
rect 12111 2150 12123 2202
rect 12175 2150 17480 2202
rect 1104 2128 17480 2150
rect 11790 2048 11796 2100
rect 11848 2088 11854 2100
rect 14090 2088 14096 2100
rect 11848 2060 14096 2088
rect 11848 2048 11854 2060
rect 14090 2048 14096 2060
rect 14148 2048 14154 2100
<< via1 >>
rect 6408 18470 6460 18522
rect 6472 18470 6524 18522
rect 6536 18470 6588 18522
rect 6600 18470 6652 18522
rect 6664 18470 6716 18522
rect 11867 18470 11919 18522
rect 11931 18470 11983 18522
rect 11995 18470 12047 18522
rect 12059 18470 12111 18522
rect 12123 18470 12175 18522
rect 2320 18300 2372 18352
rect 11612 18232 11664 18284
rect 16212 18232 16264 18284
rect 10600 18028 10652 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 15844 18028 15896 18080
rect 3679 17926 3731 17978
rect 3743 17926 3795 17978
rect 3807 17926 3859 17978
rect 3871 17926 3923 17978
rect 3935 17926 3987 17978
rect 9138 17926 9190 17978
rect 9202 17926 9254 17978
rect 9266 17926 9318 17978
rect 9330 17926 9382 17978
rect 9394 17926 9446 17978
rect 14596 17926 14648 17978
rect 14660 17926 14712 17978
rect 14724 17926 14776 17978
rect 14788 17926 14840 17978
rect 14852 17926 14904 17978
rect 6920 17824 6972 17876
rect 9588 17824 9640 17876
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 6408 17382 6460 17434
rect 6472 17382 6524 17434
rect 6536 17382 6588 17434
rect 6600 17382 6652 17434
rect 6664 17382 6716 17434
rect 11867 17382 11919 17434
rect 11931 17382 11983 17434
rect 11995 17382 12047 17434
rect 12059 17382 12111 17434
rect 12123 17382 12175 17434
rect 3679 16838 3731 16890
rect 3743 16838 3795 16890
rect 3807 16838 3859 16890
rect 3871 16838 3923 16890
rect 3935 16838 3987 16890
rect 9138 16838 9190 16890
rect 9202 16838 9254 16890
rect 9266 16838 9318 16890
rect 9330 16838 9382 16890
rect 9394 16838 9446 16890
rect 14596 16838 14648 16890
rect 14660 16838 14712 16890
rect 14724 16838 14776 16890
rect 14788 16838 14840 16890
rect 14852 16838 14904 16890
rect 6408 16294 6460 16346
rect 6472 16294 6524 16346
rect 6536 16294 6588 16346
rect 6600 16294 6652 16346
rect 6664 16294 6716 16346
rect 11867 16294 11919 16346
rect 11931 16294 11983 16346
rect 11995 16294 12047 16346
rect 12059 16294 12111 16346
rect 12123 16294 12175 16346
rect 3679 15750 3731 15802
rect 3743 15750 3795 15802
rect 3807 15750 3859 15802
rect 3871 15750 3923 15802
rect 3935 15750 3987 15802
rect 9138 15750 9190 15802
rect 9202 15750 9254 15802
rect 9266 15750 9318 15802
rect 9330 15750 9382 15802
rect 9394 15750 9446 15802
rect 14596 15750 14648 15802
rect 14660 15750 14712 15802
rect 14724 15750 14776 15802
rect 14788 15750 14840 15802
rect 14852 15750 14904 15802
rect 6408 15206 6460 15258
rect 6472 15206 6524 15258
rect 6536 15206 6588 15258
rect 6600 15206 6652 15258
rect 6664 15206 6716 15258
rect 11867 15206 11919 15258
rect 11931 15206 11983 15258
rect 11995 15206 12047 15258
rect 12059 15206 12111 15258
rect 12123 15206 12175 15258
rect 3679 14662 3731 14714
rect 3743 14662 3795 14714
rect 3807 14662 3859 14714
rect 3871 14662 3923 14714
rect 3935 14662 3987 14714
rect 9138 14662 9190 14714
rect 9202 14662 9254 14714
rect 9266 14662 9318 14714
rect 9330 14662 9382 14714
rect 9394 14662 9446 14714
rect 14596 14662 14648 14714
rect 14660 14662 14712 14714
rect 14724 14662 14776 14714
rect 14788 14662 14840 14714
rect 14852 14662 14904 14714
rect 6408 14118 6460 14170
rect 6472 14118 6524 14170
rect 6536 14118 6588 14170
rect 6600 14118 6652 14170
rect 6664 14118 6716 14170
rect 11867 14118 11919 14170
rect 11931 14118 11983 14170
rect 11995 14118 12047 14170
rect 12059 14118 12111 14170
rect 12123 14118 12175 14170
rect 3679 13574 3731 13626
rect 3743 13574 3795 13626
rect 3807 13574 3859 13626
rect 3871 13574 3923 13626
rect 3935 13574 3987 13626
rect 9138 13574 9190 13626
rect 9202 13574 9254 13626
rect 9266 13574 9318 13626
rect 9330 13574 9382 13626
rect 9394 13574 9446 13626
rect 14596 13574 14648 13626
rect 14660 13574 14712 13626
rect 14724 13574 14776 13626
rect 14788 13574 14840 13626
rect 14852 13574 14904 13626
rect 6408 13030 6460 13082
rect 6472 13030 6524 13082
rect 6536 13030 6588 13082
rect 6600 13030 6652 13082
rect 6664 13030 6716 13082
rect 11867 13030 11919 13082
rect 11931 13030 11983 13082
rect 11995 13030 12047 13082
rect 12059 13030 12111 13082
rect 12123 13030 12175 13082
rect 3679 12486 3731 12538
rect 3743 12486 3795 12538
rect 3807 12486 3859 12538
rect 3871 12486 3923 12538
rect 3935 12486 3987 12538
rect 9138 12486 9190 12538
rect 9202 12486 9254 12538
rect 9266 12486 9318 12538
rect 9330 12486 9382 12538
rect 9394 12486 9446 12538
rect 14596 12486 14648 12538
rect 14660 12486 14712 12538
rect 14724 12486 14776 12538
rect 14788 12486 14840 12538
rect 14852 12486 14904 12538
rect 6408 11942 6460 11994
rect 6472 11942 6524 11994
rect 6536 11942 6588 11994
rect 6600 11942 6652 11994
rect 6664 11942 6716 11994
rect 11867 11942 11919 11994
rect 11931 11942 11983 11994
rect 11995 11942 12047 11994
rect 12059 11942 12111 11994
rect 12123 11942 12175 11994
rect 3679 11398 3731 11450
rect 3743 11398 3795 11450
rect 3807 11398 3859 11450
rect 3871 11398 3923 11450
rect 3935 11398 3987 11450
rect 9138 11398 9190 11450
rect 9202 11398 9254 11450
rect 9266 11398 9318 11450
rect 9330 11398 9382 11450
rect 9394 11398 9446 11450
rect 14596 11398 14648 11450
rect 14660 11398 14712 11450
rect 14724 11398 14776 11450
rect 14788 11398 14840 11450
rect 14852 11398 14904 11450
rect 6408 10854 6460 10906
rect 6472 10854 6524 10906
rect 6536 10854 6588 10906
rect 6600 10854 6652 10906
rect 6664 10854 6716 10906
rect 11867 10854 11919 10906
rect 11931 10854 11983 10906
rect 11995 10854 12047 10906
rect 12059 10854 12111 10906
rect 12123 10854 12175 10906
rect 3679 10310 3731 10362
rect 3743 10310 3795 10362
rect 3807 10310 3859 10362
rect 3871 10310 3923 10362
rect 3935 10310 3987 10362
rect 9138 10310 9190 10362
rect 9202 10310 9254 10362
rect 9266 10310 9318 10362
rect 9330 10310 9382 10362
rect 9394 10310 9446 10362
rect 14596 10310 14648 10362
rect 14660 10310 14712 10362
rect 14724 10310 14776 10362
rect 14788 10310 14840 10362
rect 14852 10310 14904 10362
rect 6408 9766 6460 9818
rect 6472 9766 6524 9818
rect 6536 9766 6588 9818
rect 6600 9766 6652 9818
rect 6664 9766 6716 9818
rect 11867 9766 11919 9818
rect 11931 9766 11983 9818
rect 11995 9766 12047 9818
rect 12059 9766 12111 9818
rect 12123 9766 12175 9818
rect 3679 9222 3731 9274
rect 3743 9222 3795 9274
rect 3807 9222 3859 9274
rect 3871 9222 3923 9274
rect 3935 9222 3987 9274
rect 9138 9222 9190 9274
rect 9202 9222 9254 9274
rect 9266 9222 9318 9274
rect 9330 9222 9382 9274
rect 9394 9222 9446 9274
rect 14596 9222 14648 9274
rect 14660 9222 14712 9274
rect 14724 9222 14776 9274
rect 14788 9222 14840 9274
rect 14852 9222 14904 9274
rect 6408 8678 6460 8730
rect 6472 8678 6524 8730
rect 6536 8678 6588 8730
rect 6600 8678 6652 8730
rect 6664 8678 6716 8730
rect 11867 8678 11919 8730
rect 11931 8678 11983 8730
rect 11995 8678 12047 8730
rect 12059 8678 12111 8730
rect 12123 8678 12175 8730
rect 3679 8134 3731 8186
rect 3743 8134 3795 8186
rect 3807 8134 3859 8186
rect 3871 8134 3923 8186
rect 3935 8134 3987 8186
rect 9138 8134 9190 8186
rect 9202 8134 9254 8186
rect 9266 8134 9318 8186
rect 9330 8134 9382 8186
rect 9394 8134 9446 8186
rect 14596 8134 14648 8186
rect 14660 8134 14712 8186
rect 14724 8134 14776 8186
rect 14788 8134 14840 8186
rect 14852 8134 14904 8186
rect 6408 7590 6460 7642
rect 6472 7590 6524 7642
rect 6536 7590 6588 7642
rect 6600 7590 6652 7642
rect 6664 7590 6716 7642
rect 11867 7590 11919 7642
rect 11931 7590 11983 7642
rect 11995 7590 12047 7642
rect 12059 7590 12111 7642
rect 12123 7590 12175 7642
rect 3679 7046 3731 7098
rect 3743 7046 3795 7098
rect 3807 7046 3859 7098
rect 3871 7046 3923 7098
rect 3935 7046 3987 7098
rect 9138 7046 9190 7098
rect 9202 7046 9254 7098
rect 9266 7046 9318 7098
rect 9330 7046 9382 7098
rect 9394 7046 9446 7098
rect 14596 7046 14648 7098
rect 14660 7046 14712 7098
rect 14724 7046 14776 7098
rect 14788 7046 14840 7098
rect 14852 7046 14904 7098
rect 6408 6502 6460 6554
rect 6472 6502 6524 6554
rect 6536 6502 6588 6554
rect 6600 6502 6652 6554
rect 6664 6502 6716 6554
rect 11867 6502 11919 6554
rect 11931 6502 11983 6554
rect 11995 6502 12047 6554
rect 12059 6502 12111 6554
rect 12123 6502 12175 6554
rect 3679 5958 3731 6010
rect 3743 5958 3795 6010
rect 3807 5958 3859 6010
rect 3871 5958 3923 6010
rect 3935 5958 3987 6010
rect 9138 5958 9190 6010
rect 9202 5958 9254 6010
rect 9266 5958 9318 6010
rect 9330 5958 9382 6010
rect 9394 5958 9446 6010
rect 14596 5958 14648 6010
rect 14660 5958 14712 6010
rect 14724 5958 14776 6010
rect 14788 5958 14840 6010
rect 14852 5958 14904 6010
rect 9772 5720 9824 5772
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 11060 5652 11112 5704
rect 13084 5652 13136 5704
rect 11704 5584 11756 5636
rect 9404 5516 9456 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 11796 5516 11848 5568
rect 6408 5414 6460 5466
rect 6472 5414 6524 5466
rect 6536 5414 6588 5466
rect 6600 5414 6652 5466
rect 6664 5414 6716 5466
rect 11867 5414 11919 5466
rect 11931 5414 11983 5466
rect 11995 5414 12047 5466
rect 12059 5414 12111 5466
rect 12123 5414 12175 5466
rect 8852 5312 8904 5364
rect 9772 5312 9824 5364
rect 9404 5244 9456 5296
rect 11796 5312 11848 5364
rect 10416 5244 10468 5296
rect 11060 5176 11112 5228
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 11796 5108 11848 5160
rect 6920 4972 6972 5024
rect 3679 4870 3731 4922
rect 3743 4870 3795 4922
rect 3807 4870 3859 4922
rect 3871 4870 3923 4922
rect 3935 4870 3987 4922
rect 9138 4870 9190 4922
rect 9202 4870 9254 4922
rect 9266 4870 9318 4922
rect 9330 4870 9382 4922
rect 9394 4870 9446 4922
rect 14596 4870 14648 4922
rect 14660 4870 14712 4922
rect 14724 4870 14776 4922
rect 14788 4870 14840 4922
rect 14852 4870 14904 4922
rect 8760 4632 8812 4684
rect 7840 4564 7892 4616
rect 9588 4607 9640 4616
rect 9588 4573 9597 4607
rect 9597 4573 9631 4607
rect 9631 4573 9640 4607
rect 9588 4564 9640 4573
rect 12900 4564 12952 4616
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 15752 4564 15804 4616
rect 6736 4539 6788 4548
rect 6736 4505 6745 4539
rect 6745 4505 6779 4539
rect 6779 4505 6788 4539
rect 6736 4496 6788 4505
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 9680 4428 9732 4480
rect 14464 4471 14516 4480
rect 14464 4437 14473 4471
rect 14473 4437 14507 4471
rect 14507 4437 14516 4471
rect 14464 4428 14516 4437
rect 6408 4326 6460 4378
rect 6472 4326 6524 4378
rect 6536 4326 6588 4378
rect 6600 4326 6652 4378
rect 6664 4326 6716 4378
rect 11867 4326 11919 4378
rect 11931 4326 11983 4378
rect 11995 4326 12047 4378
rect 12059 4326 12111 4378
rect 12123 4326 12175 4378
rect 6736 4224 6788 4276
rect 7840 4267 7892 4276
rect 7840 4233 7849 4267
rect 7849 4233 7883 4267
rect 7883 4233 7892 4267
rect 7840 4224 7892 4233
rect 8484 4267 8536 4276
rect 8484 4233 8493 4267
rect 8493 4233 8527 4267
rect 8527 4233 8536 4267
rect 8484 4224 8536 4233
rect 6920 4156 6972 4208
rect 8300 4156 8352 4208
rect 7840 4088 7892 4140
rect 8024 4131 8076 4140
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 8208 4020 8260 4072
rect 8852 4088 8904 4140
rect 10600 4088 10652 4140
rect 11060 4088 11112 4140
rect 12900 4156 12952 4208
rect 14464 4156 14516 4208
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 9036 3952 9088 4004
rect 11796 4020 11848 4072
rect 12808 4063 12860 4072
rect 10232 3952 10284 4004
rect 10968 3952 11020 4004
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 6920 3884 6972 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 14924 3884 14976 3936
rect 3679 3782 3731 3834
rect 3743 3782 3795 3834
rect 3807 3782 3859 3834
rect 3871 3782 3923 3834
rect 3935 3782 3987 3834
rect 9138 3782 9190 3834
rect 9202 3782 9254 3834
rect 9266 3782 9318 3834
rect 9330 3782 9382 3834
rect 9394 3782 9446 3834
rect 14596 3782 14648 3834
rect 14660 3782 14712 3834
rect 14724 3782 14776 3834
rect 14788 3782 14840 3834
rect 14852 3782 14904 3834
rect 7840 3680 7892 3732
rect 9036 3680 9088 3732
rect 11060 3680 11112 3732
rect 12256 3680 12308 3732
rect 9680 3612 9732 3664
rect 12808 3680 12860 3732
rect 8024 3544 8076 3596
rect 12348 3544 12400 3596
rect 12440 3544 12492 3596
rect 10232 3519 10284 3528
rect 8024 3408 8076 3460
rect 8576 3408 8628 3460
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 13084 3476 13136 3528
rect 14924 3476 14976 3528
rect 11520 3408 11572 3460
rect 12532 3340 12584 3392
rect 12716 3408 12768 3460
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 12900 3340 12952 3392
rect 6408 3238 6460 3290
rect 6472 3238 6524 3290
rect 6536 3238 6588 3290
rect 6600 3238 6652 3290
rect 6664 3238 6716 3290
rect 11867 3238 11919 3290
rect 11931 3238 11983 3290
rect 11995 3238 12047 3290
rect 12059 3238 12111 3290
rect 12123 3238 12175 3290
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 7656 3068 7708 3120
rect 8392 3068 8444 3120
rect 9772 3068 9824 3120
rect 12900 3068 12952 3120
rect 8760 3000 8812 3052
rect 5724 2932 5776 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 10324 2932 10376 2984
rect 12256 2975 12308 2984
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 8760 2796 8812 2848
rect 10784 2839 10836 2848
rect 10784 2805 10793 2839
rect 10793 2805 10827 2839
rect 10827 2805 10836 2839
rect 10784 2796 10836 2805
rect 13728 2839 13780 2848
rect 13728 2805 13737 2839
rect 13737 2805 13771 2839
rect 13771 2805 13780 2839
rect 13728 2796 13780 2805
rect 3679 2694 3731 2746
rect 3743 2694 3795 2746
rect 3807 2694 3859 2746
rect 3871 2694 3923 2746
rect 3935 2694 3987 2746
rect 9138 2694 9190 2746
rect 9202 2694 9254 2746
rect 9266 2694 9318 2746
rect 9330 2694 9382 2746
rect 9394 2694 9446 2746
rect 14596 2694 14648 2746
rect 14660 2694 14712 2746
rect 14724 2694 14776 2746
rect 14788 2694 14840 2746
rect 14852 2694 14904 2746
rect 7104 2592 7156 2644
rect 8208 2592 8260 2644
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 10232 2592 10284 2644
rect 12256 2635 12308 2644
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 12532 2592 12584 2644
rect 14280 2592 14332 2644
rect 6920 2388 6972 2440
rect 1124 2320 1176 2372
rect 3424 2320 3476 2372
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 7288 2388 7340 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8576 2524 8628 2576
rect 12348 2524 12400 2576
rect 10048 2456 10100 2508
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 10784 2388 10836 2440
rect 12164 2456 12216 2508
rect 13084 2456 13136 2508
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 12808 2431 12860 2440
rect 12808 2397 12817 2431
rect 12817 2397 12851 2431
rect 12851 2397 12860 2431
rect 12808 2388 12860 2397
rect 13360 2388 13412 2440
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 9680 2320 9732 2372
rect 10416 2320 10468 2372
rect 14924 2388 14976 2440
rect 8208 2252 8260 2304
rect 10784 2252 10836 2304
rect 15016 2320 15068 2372
rect 13728 2252 13780 2304
rect 17316 2320 17368 2372
rect 6408 2150 6460 2202
rect 6472 2150 6524 2202
rect 6536 2150 6588 2202
rect 6600 2150 6652 2202
rect 6664 2150 6716 2202
rect 11867 2150 11919 2202
rect 11931 2150 11983 2202
rect 11995 2150 12047 2202
rect 12059 2150 12111 2202
rect 12123 2150 12175 2202
rect 11796 2048 11848 2100
rect 14096 2048 14148 2100
<< metal2 >>
rect 2318 19931 2374 20731
rect 6918 19931 6974 20731
rect 11610 19931 11666 20731
rect 16210 19931 16266 20731
rect 2332 18358 2360 19931
rect 6408 18524 6716 18544
rect 6408 18522 6414 18524
rect 6470 18522 6494 18524
rect 6550 18522 6574 18524
rect 6630 18522 6654 18524
rect 6710 18522 6716 18524
rect 6470 18470 6472 18522
rect 6652 18470 6654 18522
rect 6408 18468 6414 18470
rect 6470 18468 6494 18470
rect 6550 18468 6574 18470
rect 6630 18468 6654 18470
rect 6710 18468 6716 18470
rect 6408 18448 6716 18468
rect 2320 18352 2372 18358
rect 2320 18294 2372 18300
rect 3679 17980 3987 18000
rect 3679 17978 3685 17980
rect 3741 17978 3765 17980
rect 3821 17978 3845 17980
rect 3901 17978 3925 17980
rect 3981 17978 3987 17980
rect 3741 17926 3743 17978
rect 3923 17926 3925 17978
rect 3679 17924 3685 17926
rect 3741 17924 3765 17926
rect 3821 17924 3845 17926
rect 3901 17924 3925 17926
rect 3981 17924 3987 17926
rect 3679 17904 3987 17924
rect 6932 17882 6960 19931
rect 11624 18290 11652 19931
rect 11867 18524 12175 18544
rect 11867 18522 11873 18524
rect 11929 18522 11953 18524
rect 12009 18522 12033 18524
rect 12089 18522 12113 18524
rect 12169 18522 12175 18524
rect 11929 18470 11931 18522
rect 12111 18470 12113 18522
rect 11867 18468 11873 18470
rect 11929 18468 11953 18470
rect 12009 18468 12033 18470
rect 12089 18468 12113 18470
rect 12169 18468 12175 18470
rect 11867 18448 12175 18468
rect 16224 18290 16252 19931
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 9138 17980 9446 18000
rect 9138 17978 9144 17980
rect 9200 17978 9224 17980
rect 9280 17978 9304 17980
rect 9360 17978 9384 17980
rect 9440 17978 9446 17980
rect 9200 17926 9202 17978
rect 9382 17926 9384 17978
rect 9138 17924 9144 17926
rect 9200 17924 9224 17926
rect 9280 17924 9304 17926
rect 9360 17924 9384 17926
rect 9440 17924 9446 17926
rect 9138 17904 9446 17924
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 6408 17436 6716 17456
rect 6408 17434 6414 17436
rect 6470 17434 6494 17436
rect 6550 17434 6574 17436
rect 6630 17434 6654 17436
rect 6710 17434 6716 17436
rect 6470 17382 6472 17434
rect 6652 17382 6654 17434
rect 6408 17380 6414 17382
rect 6470 17380 6494 17382
rect 6550 17380 6574 17382
rect 6630 17380 6654 17382
rect 6710 17380 6716 17382
rect 6408 17360 6716 17380
rect 3679 16892 3987 16912
rect 3679 16890 3685 16892
rect 3741 16890 3765 16892
rect 3821 16890 3845 16892
rect 3901 16890 3925 16892
rect 3981 16890 3987 16892
rect 3741 16838 3743 16890
rect 3923 16838 3925 16890
rect 3679 16836 3685 16838
rect 3741 16836 3765 16838
rect 3821 16836 3845 16838
rect 3901 16836 3925 16838
rect 3981 16836 3987 16838
rect 3679 16816 3987 16836
rect 9138 16892 9446 16912
rect 9138 16890 9144 16892
rect 9200 16890 9224 16892
rect 9280 16890 9304 16892
rect 9360 16890 9384 16892
rect 9440 16890 9446 16892
rect 9200 16838 9202 16890
rect 9382 16838 9384 16890
rect 9138 16836 9144 16838
rect 9200 16836 9224 16838
rect 9280 16836 9304 16838
rect 9360 16836 9384 16838
rect 9440 16836 9446 16838
rect 9138 16816 9446 16836
rect 6408 16348 6716 16368
rect 6408 16346 6414 16348
rect 6470 16346 6494 16348
rect 6550 16346 6574 16348
rect 6630 16346 6654 16348
rect 6710 16346 6716 16348
rect 6470 16294 6472 16346
rect 6652 16294 6654 16346
rect 6408 16292 6414 16294
rect 6470 16292 6494 16294
rect 6550 16292 6574 16294
rect 6630 16292 6654 16294
rect 6710 16292 6716 16294
rect 6408 16272 6716 16292
rect 3679 15804 3987 15824
rect 3679 15802 3685 15804
rect 3741 15802 3765 15804
rect 3821 15802 3845 15804
rect 3901 15802 3925 15804
rect 3981 15802 3987 15804
rect 3741 15750 3743 15802
rect 3923 15750 3925 15802
rect 3679 15748 3685 15750
rect 3741 15748 3765 15750
rect 3821 15748 3845 15750
rect 3901 15748 3925 15750
rect 3981 15748 3987 15750
rect 3679 15728 3987 15748
rect 9138 15804 9446 15824
rect 9138 15802 9144 15804
rect 9200 15802 9224 15804
rect 9280 15802 9304 15804
rect 9360 15802 9384 15804
rect 9440 15802 9446 15804
rect 9200 15750 9202 15802
rect 9382 15750 9384 15802
rect 9138 15748 9144 15750
rect 9200 15748 9224 15750
rect 9280 15748 9304 15750
rect 9360 15748 9384 15750
rect 9440 15748 9446 15750
rect 9138 15728 9446 15748
rect 6408 15260 6716 15280
rect 6408 15258 6414 15260
rect 6470 15258 6494 15260
rect 6550 15258 6574 15260
rect 6630 15258 6654 15260
rect 6710 15258 6716 15260
rect 6470 15206 6472 15258
rect 6652 15206 6654 15258
rect 6408 15204 6414 15206
rect 6470 15204 6494 15206
rect 6550 15204 6574 15206
rect 6630 15204 6654 15206
rect 6710 15204 6716 15206
rect 6408 15184 6716 15204
rect 3679 14716 3987 14736
rect 3679 14714 3685 14716
rect 3741 14714 3765 14716
rect 3821 14714 3845 14716
rect 3901 14714 3925 14716
rect 3981 14714 3987 14716
rect 3741 14662 3743 14714
rect 3923 14662 3925 14714
rect 3679 14660 3685 14662
rect 3741 14660 3765 14662
rect 3821 14660 3845 14662
rect 3901 14660 3925 14662
rect 3981 14660 3987 14662
rect 3679 14640 3987 14660
rect 9138 14716 9446 14736
rect 9138 14714 9144 14716
rect 9200 14714 9224 14716
rect 9280 14714 9304 14716
rect 9360 14714 9384 14716
rect 9440 14714 9446 14716
rect 9200 14662 9202 14714
rect 9382 14662 9384 14714
rect 9138 14660 9144 14662
rect 9200 14660 9224 14662
rect 9280 14660 9304 14662
rect 9360 14660 9384 14662
rect 9440 14660 9446 14662
rect 9138 14640 9446 14660
rect 6408 14172 6716 14192
rect 6408 14170 6414 14172
rect 6470 14170 6494 14172
rect 6550 14170 6574 14172
rect 6630 14170 6654 14172
rect 6710 14170 6716 14172
rect 6470 14118 6472 14170
rect 6652 14118 6654 14170
rect 6408 14116 6414 14118
rect 6470 14116 6494 14118
rect 6550 14116 6574 14118
rect 6630 14116 6654 14118
rect 6710 14116 6716 14118
rect 6408 14096 6716 14116
rect 3679 13628 3987 13648
rect 3679 13626 3685 13628
rect 3741 13626 3765 13628
rect 3821 13626 3845 13628
rect 3901 13626 3925 13628
rect 3981 13626 3987 13628
rect 3741 13574 3743 13626
rect 3923 13574 3925 13626
rect 3679 13572 3685 13574
rect 3741 13572 3765 13574
rect 3821 13572 3845 13574
rect 3901 13572 3925 13574
rect 3981 13572 3987 13574
rect 3679 13552 3987 13572
rect 9138 13628 9446 13648
rect 9138 13626 9144 13628
rect 9200 13626 9224 13628
rect 9280 13626 9304 13628
rect 9360 13626 9384 13628
rect 9440 13626 9446 13628
rect 9200 13574 9202 13626
rect 9382 13574 9384 13626
rect 9138 13572 9144 13574
rect 9200 13572 9224 13574
rect 9280 13572 9304 13574
rect 9360 13572 9384 13574
rect 9440 13572 9446 13574
rect 9138 13552 9446 13572
rect 6408 13084 6716 13104
rect 6408 13082 6414 13084
rect 6470 13082 6494 13084
rect 6550 13082 6574 13084
rect 6630 13082 6654 13084
rect 6710 13082 6716 13084
rect 6470 13030 6472 13082
rect 6652 13030 6654 13082
rect 6408 13028 6414 13030
rect 6470 13028 6494 13030
rect 6550 13028 6574 13030
rect 6630 13028 6654 13030
rect 6710 13028 6716 13030
rect 6408 13008 6716 13028
rect 3679 12540 3987 12560
rect 3679 12538 3685 12540
rect 3741 12538 3765 12540
rect 3821 12538 3845 12540
rect 3901 12538 3925 12540
rect 3981 12538 3987 12540
rect 3741 12486 3743 12538
rect 3923 12486 3925 12538
rect 3679 12484 3685 12486
rect 3741 12484 3765 12486
rect 3821 12484 3845 12486
rect 3901 12484 3925 12486
rect 3981 12484 3987 12486
rect 3679 12464 3987 12484
rect 9138 12540 9446 12560
rect 9138 12538 9144 12540
rect 9200 12538 9224 12540
rect 9280 12538 9304 12540
rect 9360 12538 9384 12540
rect 9440 12538 9446 12540
rect 9200 12486 9202 12538
rect 9382 12486 9384 12538
rect 9138 12484 9144 12486
rect 9200 12484 9224 12486
rect 9280 12484 9304 12486
rect 9360 12484 9384 12486
rect 9440 12484 9446 12486
rect 9138 12464 9446 12484
rect 6408 11996 6716 12016
rect 6408 11994 6414 11996
rect 6470 11994 6494 11996
rect 6550 11994 6574 11996
rect 6630 11994 6654 11996
rect 6710 11994 6716 11996
rect 6470 11942 6472 11994
rect 6652 11942 6654 11994
rect 6408 11940 6414 11942
rect 6470 11940 6494 11942
rect 6550 11940 6574 11942
rect 6630 11940 6654 11942
rect 6710 11940 6716 11942
rect 6408 11920 6716 11940
rect 3679 11452 3987 11472
rect 3679 11450 3685 11452
rect 3741 11450 3765 11452
rect 3821 11450 3845 11452
rect 3901 11450 3925 11452
rect 3981 11450 3987 11452
rect 3741 11398 3743 11450
rect 3923 11398 3925 11450
rect 3679 11396 3685 11398
rect 3741 11396 3765 11398
rect 3821 11396 3845 11398
rect 3901 11396 3925 11398
rect 3981 11396 3987 11398
rect 3679 11376 3987 11396
rect 9138 11452 9446 11472
rect 9138 11450 9144 11452
rect 9200 11450 9224 11452
rect 9280 11450 9304 11452
rect 9360 11450 9384 11452
rect 9440 11450 9446 11452
rect 9200 11398 9202 11450
rect 9382 11398 9384 11450
rect 9138 11396 9144 11398
rect 9200 11396 9224 11398
rect 9280 11396 9304 11398
rect 9360 11396 9384 11398
rect 9440 11396 9446 11398
rect 9138 11376 9446 11396
rect 6408 10908 6716 10928
rect 6408 10906 6414 10908
rect 6470 10906 6494 10908
rect 6550 10906 6574 10908
rect 6630 10906 6654 10908
rect 6710 10906 6716 10908
rect 6470 10854 6472 10906
rect 6652 10854 6654 10906
rect 6408 10852 6414 10854
rect 6470 10852 6494 10854
rect 6550 10852 6574 10854
rect 6630 10852 6654 10854
rect 6710 10852 6716 10854
rect 6408 10832 6716 10852
rect 3679 10364 3987 10384
rect 3679 10362 3685 10364
rect 3741 10362 3765 10364
rect 3821 10362 3845 10364
rect 3901 10362 3925 10364
rect 3981 10362 3987 10364
rect 3741 10310 3743 10362
rect 3923 10310 3925 10362
rect 3679 10308 3685 10310
rect 3741 10308 3765 10310
rect 3821 10308 3845 10310
rect 3901 10308 3925 10310
rect 3981 10308 3987 10310
rect 3679 10288 3987 10308
rect 9138 10364 9446 10384
rect 9138 10362 9144 10364
rect 9200 10362 9224 10364
rect 9280 10362 9304 10364
rect 9360 10362 9384 10364
rect 9440 10362 9446 10364
rect 9200 10310 9202 10362
rect 9382 10310 9384 10362
rect 9138 10308 9144 10310
rect 9200 10308 9224 10310
rect 9280 10308 9304 10310
rect 9360 10308 9384 10310
rect 9440 10308 9446 10310
rect 9138 10288 9446 10308
rect 6408 9820 6716 9840
rect 6408 9818 6414 9820
rect 6470 9818 6494 9820
rect 6550 9818 6574 9820
rect 6630 9818 6654 9820
rect 6710 9818 6716 9820
rect 6470 9766 6472 9818
rect 6652 9766 6654 9818
rect 6408 9764 6414 9766
rect 6470 9764 6494 9766
rect 6550 9764 6574 9766
rect 6630 9764 6654 9766
rect 6710 9764 6716 9766
rect 6408 9744 6716 9764
rect 3679 9276 3987 9296
rect 3679 9274 3685 9276
rect 3741 9274 3765 9276
rect 3821 9274 3845 9276
rect 3901 9274 3925 9276
rect 3981 9274 3987 9276
rect 3741 9222 3743 9274
rect 3923 9222 3925 9274
rect 3679 9220 3685 9222
rect 3741 9220 3765 9222
rect 3821 9220 3845 9222
rect 3901 9220 3925 9222
rect 3981 9220 3987 9222
rect 3679 9200 3987 9220
rect 9138 9276 9446 9296
rect 9138 9274 9144 9276
rect 9200 9274 9224 9276
rect 9280 9274 9304 9276
rect 9360 9274 9384 9276
rect 9440 9274 9446 9276
rect 9200 9222 9202 9274
rect 9382 9222 9384 9274
rect 9138 9220 9144 9222
rect 9200 9220 9224 9222
rect 9280 9220 9304 9222
rect 9360 9220 9384 9222
rect 9440 9220 9446 9222
rect 9138 9200 9446 9220
rect 6408 8732 6716 8752
rect 6408 8730 6414 8732
rect 6470 8730 6494 8732
rect 6550 8730 6574 8732
rect 6630 8730 6654 8732
rect 6710 8730 6716 8732
rect 6470 8678 6472 8730
rect 6652 8678 6654 8730
rect 6408 8676 6414 8678
rect 6470 8676 6494 8678
rect 6550 8676 6574 8678
rect 6630 8676 6654 8678
rect 6710 8676 6716 8678
rect 6408 8656 6716 8676
rect 3679 8188 3987 8208
rect 3679 8186 3685 8188
rect 3741 8186 3765 8188
rect 3821 8186 3845 8188
rect 3901 8186 3925 8188
rect 3981 8186 3987 8188
rect 3741 8134 3743 8186
rect 3923 8134 3925 8186
rect 3679 8132 3685 8134
rect 3741 8132 3765 8134
rect 3821 8132 3845 8134
rect 3901 8132 3925 8134
rect 3981 8132 3987 8134
rect 3679 8112 3987 8132
rect 9138 8188 9446 8208
rect 9138 8186 9144 8188
rect 9200 8186 9224 8188
rect 9280 8186 9304 8188
rect 9360 8186 9384 8188
rect 9440 8186 9446 8188
rect 9200 8134 9202 8186
rect 9382 8134 9384 8186
rect 9138 8132 9144 8134
rect 9200 8132 9224 8134
rect 9280 8132 9304 8134
rect 9360 8132 9384 8134
rect 9440 8132 9446 8134
rect 9138 8112 9446 8132
rect 6408 7644 6716 7664
rect 6408 7642 6414 7644
rect 6470 7642 6494 7644
rect 6550 7642 6574 7644
rect 6630 7642 6654 7644
rect 6710 7642 6716 7644
rect 6470 7590 6472 7642
rect 6652 7590 6654 7642
rect 6408 7588 6414 7590
rect 6470 7588 6494 7590
rect 6550 7588 6574 7590
rect 6630 7588 6654 7590
rect 6710 7588 6716 7590
rect 6408 7568 6716 7588
rect 3679 7100 3987 7120
rect 3679 7098 3685 7100
rect 3741 7098 3765 7100
rect 3821 7098 3845 7100
rect 3901 7098 3925 7100
rect 3981 7098 3987 7100
rect 3741 7046 3743 7098
rect 3923 7046 3925 7098
rect 3679 7044 3685 7046
rect 3741 7044 3765 7046
rect 3821 7044 3845 7046
rect 3901 7044 3925 7046
rect 3981 7044 3987 7046
rect 3679 7024 3987 7044
rect 9138 7100 9446 7120
rect 9138 7098 9144 7100
rect 9200 7098 9224 7100
rect 9280 7098 9304 7100
rect 9360 7098 9384 7100
rect 9440 7098 9446 7100
rect 9200 7046 9202 7098
rect 9382 7046 9384 7098
rect 9138 7044 9144 7046
rect 9200 7044 9224 7046
rect 9280 7044 9304 7046
rect 9360 7044 9384 7046
rect 9440 7044 9446 7046
rect 9138 7024 9446 7044
rect 6408 6556 6716 6576
rect 6408 6554 6414 6556
rect 6470 6554 6494 6556
rect 6550 6554 6574 6556
rect 6630 6554 6654 6556
rect 6710 6554 6716 6556
rect 6470 6502 6472 6554
rect 6652 6502 6654 6554
rect 6408 6500 6414 6502
rect 6470 6500 6494 6502
rect 6550 6500 6574 6502
rect 6630 6500 6654 6502
rect 6710 6500 6716 6502
rect 6408 6480 6716 6500
rect 3679 6012 3987 6032
rect 3679 6010 3685 6012
rect 3741 6010 3765 6012
rect 3821 6010 3845 6012
rect 3901 6010 3925 6012
rect 3981 6010 3987 6012
rect 3741 5958 3743 6010
rect 3923 5958 3925 6010
rect 3679 5956 3685 5958
rect 3741 5956 3765 5958
rect 3821 5956 3845 5958
rect 3901 5956 3925 5958
rect 3981 5956 3987 5958
rect 3679 5936 3987 5956
rect 9138 6012 9446 6032
rect 9138 6010 9144 6012
rect 9200 6010 9224 6012
rect 9280 6010 9304 6012
rect 9360 6010 9384 6012
rect 9440 6010 9446 6012
rect 9200 5958 9202 6010
rect 9382 5958 9384 6010
rect 9138 5956 9144 5958
rect 9200 5956 9224 5958
rect 9280 5956 9304 5958
rect 9360 5956 9384 5958
rect 9440 5956 9446 5958
rect 9138 5936 9446 5956
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 6408 5468 6716 5488
rect 6408 5466 6414 5468
rect 6470 5466 6494 5468
rect 6550 5466 6574 5468
rect 6630 5466 6654 5468
rect 6710 5466 6716 5468
rect 6470 5414 6472 5466
rect 6652 5414 6654 5466
rect 6408 5412 6414 5414
rect 6470 5412 6494 5414
rect 6550 5412 6574 5414
rect 6630 5412 6654 5414
rect 6710 5412 6716 5414
rect 6408 5392 6716 5412
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 3679 4924 3987 4944
rect 3679 4922 3685 4924
rect 3741 4922 3765 4924
rect 3821 4922 3845 4924
rect 3901 4922 3925 4924
rect 3981 4922 3987 4924
rect 3741 4870 3743 4922
rect 3923 4870 3925 4922
rect 3679 4868 3685 4870
rect 3741 4868 3765 4870
rect 3821 4868 3845 4870
rect 3901 4868 3925 4870
rect 3981 4868 3987 4870
rect 3679 4848 3987 4868
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6408 4380 6716 4400
rect 6408 4378 6414 4380
rect 6470 4378 6494 4380
rect 6550 4378 6574 4380
rect 6630 4378 6654 4380
rect 6710 4378 6716 4380
rect 6470 4326 6472 4378
rect 6652 4326 6654 4378
rect 6408 4324 6414 4326
rect 6470 4324 6494 4326
rect 6550 4324 6574 4326
rect 6630 4324 6654 4326
rect 6710 4324 6716 4326
rect 6408 4304 6716 4324
rect 6748 4282 6776 4490
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6932 4214 6960 4966
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 4282 7880 4558
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6932 3942 6960 4150
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 3679 3836 3987 3856
rect 3679 3834 3685 3836
rect 3741 3834 3765 3836
rect 3821 3834 3845 3836
rect 3901 3834 3925 3836
rect 3981 3834 3987 3836
rect 3741 3782 3743 3834
rect 3923 3782 3925 3834
rect 3679 3780 3685 3782
rect 3741 3780 3765 3782
rect 3821 3780 3845 3782
rect 3901 3780 3925 3782
rect 3981 3780 3987 3782
rect 3679 3760 3987 3780
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 2990 5764 3334
rect 6408 3292 6716 3312
rect 6408 3290 6414 3292
rect 6470 3290 6494 3292
rect 6550 3290 6574 3292
rect 6630 3290 6654 3292
rect 6710 3290 6716 3292
rect 6470 3238 6472 3290
rect 6652 3238 6654 3290
rect 6408 3236 6414 3238
rect 6470 3236 6494 3238
rect 6550 3236 6574 3238
rect 6630 3236 6654 3238
rect 6710 3236 6716 3238
rect 6408 3216 6716 3236
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 3679 2748 3987 2768
rect 3679 2746 3685 2748
rect 3741 2746 3765 2748
rect 3821 2746 3845 2748
rect 3901 2746 3925 2748
rect 3981 2746 3987 2748
rect 3741 2694 3743 2746
rect 3923 2694 3925 2746
rect 3679 2692 3685 2694
rect 3741 2692 3765 2694
rect 3821 2692 3845 2694
rect 3901 2692 3925 2694
rect 3981 2692 3987 2694
rect 3679 2672 3987 2692
rect 6932 2446 6960 3878
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7116 2650 7144 2926
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7300 2446 7328 4014
rect 7852 3738 7880 4082
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 3126 7696 3334
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7852 2446 7880 3674
rect 8036 3602 8064 4082
rect 8220 4078 8248 4422
rect 8496 4282 8524 5102
rect 8772 4690 8800 5102
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 1124 2372 1176 2378
rect 1124 2314 1176 2320
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 1136 800 1164 2314
rect 3436 800 3464 2314
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5644 1170 5672 2246
rect 6408 2204 6716 2224
rect 6408 2202 6414 2204
rect 6470 2202 6494 2204
rect 6550 2202 6574 2204
rect 6630 2202 6654 2204
rect 6710 2202 6716 2204
rect 6470 2150 6472 2202
rect 6652 2150 6654 2202
rect 6408 2148 6414 2150
rect 6470 2148 6494 2150
rect 6550 2148 6574 2150
rect 6630 2148 6654 2150
rect 6710 2148 6716 2150
rect 6408 2128 6716 2148
rect 5644 1142 5764 1170
rect 5736 800 5764 1142
rect 8036 800 8064 3402
rect 8312 2666 8340 4150
rect 8576 3460 8628 3466
rect 8576 3402 8628 3408
rect 8588 3194 8616 3402
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8220 2650 8340 2666
rect 8404 2650 8432 3062
rect 8208 2644 8340 2650
rect 8260 2638 8340 2644
rect 8392 2644 8444 2650
rect 8208 2586 8260 2592
rect 8392 2586 8444 2592
rect 8588 2582 8616 3130
rect 8772 3058 8800 4626
rect 8864 4146 8892 5306
rect 9416 5302 9444 5510
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9138 4924 9446 4944
rect 9138 4922 9144 4924
rect 9200 4922 9224 4924
rect 9280 4922 9304 4924
rect 9360 4922 9384 4924
rect 9440 4922 9446 4924
rect 9200 4870 9202 4922
rect 9382 4870 9384 4922
rect 9138 4868 9144 4870
rect 9200 4868 9224 4870
rect 9280 4868 9304 4870
rect 9360 4868 9384 4870
rect 9440 4868 9446 4870
rect 9138 4848 9446 4868
rect 9600 4622 9628 17818
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9784 5370 9812 5714
rect 10612 5710 10640 18022
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 10428 5302 10456 5510
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 9048 3738 9076 3946
rect 9138 3836 9446 3856
rect 9138 3834 9144 3836
rect 9200 3834 9224 3836
rect 9280 3834 9304 3836
rect 9360 3834 9384 3836
rect 9440 3834 9446 3836
rect 9200 3782 9202 3834
rect 9382 3782 9384 3834
rect 9138 3780 9144 3782
rect 9200 3780 9224 3782
rect 9280 3780 9304 3782
rect 9360 3780 9384 3782
rect 9440 3780 9446 3782
rect 9138 3760 9446 3780
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9692 3670 9720 4422
rect 10612 4146 10640 5646
rect 11072 5234 11100 5646
rect 11716 5642 11744 18022
rect 14596 17980 14904 18000
rect 14596 17978 14602 17980
rect 14658 17978 14682 17980
rect 14738 17978 14762 17980
rect 14818 17978 14842 17980
rect 14898 17978 14904 17980
rect 14658 17926 14660 17978
rect 14840 17926 14842 17978
rect 14596 17924 14602 17926
rect 14658 17924 14682 17926
rect 14738 17924 14762 17926
rect 14818 17924 14842 17926
rect 14898 17924 14904 17926
rect 14596 17904 14904 17924
rect 15856 17678 15884 18022
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 11867 17436 12175 17456
rect 11867 17434 11873 17436
rect 11929 17434 11953 17436
rect 12009 17434 12033 17436
rect 12089 17434 12113 17436
rect 12169 17434 12175 17436
rect 11929 17382 11931 17434
rect 12111 17382 12113 17434
rect 11867 17380 11873 17382
rect 11929 17380 11953 17382
rect 12009 17380 12033 17382
rect 12089 17380 12113 17382
rect 12169 17380 12175 17382
rect 11867 17360 12175 17380
rect 14596 16892 14904 16912
rect 14596 16890 14602 16892
rect 14658 16890 14682 16892
rect 14738 16890 14762 16892
rect 14818 16890 14842 16892
rect 14898 16890 14904 16892
rect 14658 16838 14660 16890
rect 14840 16838 14842 16890
rect 14596 16836 14602 16838
rect 14658 16836 14682 16838
rect 14738 16836 14762 16838
rect 14818 16836 14842 16838
rect 14898 16836 14904 16838
rect 14596 16816 14904 16836
rect 11867 16348 12175 16368
rect 11867 16346 11873 16348
rect 11929 16346 11953 16348
rect 12009 16346 12033 16348
rect 12089 16346 12113 16348
rect 12169 16346 12175 16348
rect 11929 16294 11931 16346
rect 12111 16294 12113 16346
rect 11867 16292 11873 16294
rect 11929 16292 11953 16294
rect 12009 16292 12033 16294
rect 12089 16292 12113 16294
rect 12169 16292 12175 16294
rect 11867 16272 12175 16292
rect 14596 15804 14904 15824
rect 14596 15802 14602 15804
rect 14658 15802 14682 15804
rect 14738 15802 14762 15804
rect 14818 15802 14842 15804
rect 14898 15802 14904 15804
rect 14658 15750 14660 15802
rect 14840 15750 14842 15802
rect 14596 15748 14602 15750
rect 14658 15748 14682 15750
rect 14738 15748 14762 15750
rect 14818 15748 14842 15750
rect 14898 15748 14904 15750
rect 14596 15728 14904 15748
rect 11867 15260 12175 15280
rect 11867 15258 11873 15260
rect 11929 15258 11953 15260
rect 12009 15258 12033 15260
rect 12089 15258 12113 15260
rect 12169 15258 12175 15260
rect 11929 15206 11931 15258
rect 12111 15206 12113 15258
rect 11867 15204 11873 15206
rect 11929 15204 11953 15206
rect 12009 15204 12033 15206
rect 12089 15204 12113 15206
rect 12169 15204 12175 15206
rect 11867 15184 12175 15204
rect 14596 14716 14904 14736
rect 14596 14714 14602 14716
rect 14658 14714 14682 14716
rect 14738 14714 14762 14716
rect 14818 14714 14842 14716
rect 14898 14714 14904 14716
rect 14658 14662 14660 14714
rect 14840 14662 14842 14714
rect 14596 14660 14602 14662
rect 14658 14660 14682 14662
rect 14738 14660 14762 14662
rect 14818 14660 14842 14662
rect 14898 14660 14904 14662
rect 14596 14640 14904 14660
rect 11867 14172 12175 14192
rect 11867 14170 11873 14172
rect 11929 14170 11953 14172
rect 12009 14170 12033 14172
rect 12089 14170 12113 14172
rect 12169 14170 12175 14172
rect 11929 14118 11931 14170
rect 12111 14118 12113 14170
rect 11867 14116 11873 14118
rect 11929 14116 11953 14118
rect 12009 14116 12033 14118
rect 12089 14116 12113 14118
rect 12169 14116 12175 14118
rect 11867 14096 12175 14116
rect 14596 13628 14904 13648
rect 14596 13626 14602 13628
rect 14658 13626 14682 13628
rect 14738 13626 14762 13628
rect 14818 13626 14842 13628
rect 14898 13626 14904 13628
rect 14658 13574 14660 13626
rect 14840 13574 14842 13626
rect 14596 13572 14602 13574
rect 14658 13572 14682 13574
rect 14738 13572 14762 13574
rect 14818 13572 14842 13574
rect 14898 13572 14904 13574
rect 14596 13552 14904 13572
rect 11867 13084 12175 13104
rect 11867 13082 11873 13084
rect 11929 13082 11953 13084
rect 12009 13082 12033 13084
rect 12089 13082 12113 13084
rect 12169 13082 12175 13084
rect 11929 13030 11931 13082
rect 12111 13030 12113 13082
rect 11867 13028 11873 13030
rect 11929 13028 11953 13030
rect 12009 13028 12033 13030
rect 12089 13028 12113 13030
rect 12169 13028 12175 13030
rect 11867 13008 12175 13028
rect 14596 12540 14904 12560
rect 14596 12538 14602 12540
rect 14658 12538 14682 12540
rect 14738 12538 14762 12540
rect 14818 12538 14842 12540
rect 14898 12538 14904 12540
rect 14658 12486 14660 12538
rect 14840 12486 14842 12538
rect 14596 12484 14602 12486
rect 14658 12484 14682 12486
rect 14738 12484 14762 12486
rect 14818 12484 14842 12486
rect 14898 12484 14904 12486
rect 14596 12464 14904 12484
rect 11867 11996 12175 12016
rect 11867 11994 11873 11996
rect 11929 11994 11953 11996
rect 12009 11994 12033 11996
rect 12089 11994 12113 11996
rect 12169 11994 12175 11996
rect 11929 11942 11931 11994
rect 12111 11942 12113 11994
rect 11867 11940 11873 11942
rect 11929 11940 11953 11942
rect 12009 11940 12033 11942
rect 12089 11940 12113 11942
rect 12169 11940 12175 11942
rect 11867 11920 12175 11940
rect 14596 11452 14904 11472
rect 14596 11450 14602 11452
rect 14658 11450 14682 11452
rect 14738 11450 14762 11452
rect 14818 11450 14842 11452
rect 14898 11450 14904 11452
rect 14658 11398 14660 11450
rect 14840 11398 14842 11450
rect 14596 11396 14602 11398
rect 14658 11396 14682 11398
rect 14738 11396 14762 11398
rect 14818 11396 14842 11398
rect 14898 11396 14904 11398
rect 14596 11376 14904 11396
rect 11867 10908 12175 10928
rect 11867 10906 11873 10908
rect 11929 10906 11953 10908
rect 12009 10906 12033 10908
rect 12089 10906 12113 10908
rect 12169 10906 12175 10908
rect 11929 10854 11931 10906
rect 12111 10854 12113 10906
rect 11867 10852 11873 10854
rect 11929 10852 11953 10854
rect 12009 10852 12033 10854
rect 12089 10852 12113 10854
rect 12169 10852 12175 10854
rect 11867 10832 12175 10852
rect 14596 10364 14904 10384
rect 14596 10362 14602 10364
rect 14658 10362 14682 10364
rect 14738 10362 14762 10364
rect 14818 10362 14842 10364
rect 14898 10362 14904 10364
rect 14658 10310 14660 10362
rect 14840 10310 14842 10362
rect 14596 10308 14602 10310
rect 14658 10308 14682 10310
rect 14738 10308 14762 10310
rect 14818 10308 14842 10310
rect 14898 10308 14904 10310
rect 14596 10288 14904 10308
rect 11867 9820 12175 9840
rect 11867 9818 11873 9820
rect 11929 9818 11953 9820
rect 12009 9818 12033 9820
rect 12089 9818 12113 9820
rect 12169 9818 12175 9820
rect 11929 9766 11931 9818
rect 12111 9766 12113 9818
rect 11867 9764 11873 9766
rect 11929 9764 11953 9766
rect 12009 9764 12033 9766
rect 12089 9764 12113 9766
rect 12169 9764 12175 9766
rect 11867 9744 12175 9764
rect 14596 9276 14904 9296
rect 14596 9274 14602 9276
rect 14658 9274 14682 9276
rect 14738 9274 14762 9276
rect 14818 9274 14842 9276
rect 14898 9274 14904 9276
rect 14658 9222 14660 9274
rect 14840 9222 14842 9274
rect 14596 9220 14602 9222
rect 14658 9220 14682 9222
rect 14738 9220 14762 9222
rect 14818 9220 14842 9222
rect 14898 9220 14904 9222
rect 14596 9200 14904 9220
rect 11867 8732 12175 8752
rect 11867 8730 11873 8732
rect 11929 8730 11953 8732
rect 12009 8730 12033 8732
rect 12089 8730 12113 8732
rect 12169 8730 12175 8732
rect 11929 8678 11931 8730
rect 12111 8678 12113 8730
rect 11867 8676 11873 8678
rect 11929 8676 11953 8678
rect 12009 8676 12033 8678
rect 12089 8676 12113 8678
rect 12169 8676 12175 8678
rect 11867 8656 12175 8676
rect 14596 8188 14904 8208
rect 14596 8186 14602 8188
rect 14658 8186 14682 8188
rect 14738 8186 14762 8188
rect 14818 8186 14842 8188
rect 14898 8186 14904 8188
rect 14658 8134 14660 8186
rect 14840 8134 14842 8186
rect 14596 8132 14602 8134
rect 14658 8132 14682 8134
rect 14738 8132 14762 8134
rect 14818 8132 14842 8134
rect 14898 8132 14904 8134
rect 14596 8112 14904 8132
rect 11867 7644 12175 7664
rect 11867 7642 11873 7644
rect 11929 7642 11953 7644
rect 12009 7642 12033 7644
rect 12089 7642 12113 7644
rect 12169 7642 12175 7644
rect 11929 7590 11931 7642
rect 12111 7590 12113 7642
rect 11867 7588 11873 7590
rect 11929 7588 11953 7590
rect 12009 7588 12033 7590
rect 12089 7588 12113 7590
rect 12169 7588 12175 7590
rect 11867 7568 12175 7588
rect 14596 7100 14904 7120
rect 14596 7098 14602 7100
rect 14658 7098 14682 7100
rect 14738 7098 14762 7100
rect 14818 7098 14842 7100
rect 14898 7098 14904 7100
rect 14658 7046 14660 7098
rect 14840 7046 14842 7098
rect 14596 7044 14602 7046
rect 14658 7044 14682 7046
rect 14738 7044 14762 7046
rect 14818 7044 14842 7046
rect 14898 7044 14904 7046
rect 14596 7024 14904 7044
rect 11867 6556 12175 6576
rect 11867 6554 11873 6556
rect 11929 6554 11953 6556
rect 12009 6554 12033 6556
rect 12089 6554 12113 6556
rect 12169 6554 12175 6556
rect 11929 6502 11931 6554
rect 12111 6502 12113 6554
rect 11867 6500 11873 6502
rect 11929 6500 11953 6502
rect 12009 6500 12033 6502
rect 12089 6500 12113 6502
rect 12169 6500 12175 6502
rect 11867 6480 12175 6500
rect 14596 6012 14904 6032
rect 14596 6010 14602 6012
rect 14658 6010 14682 6012
rect 14738 6010 14762 6012
rect 14818 6010 14842 6012
rect 14898 6010 14904 6012
rect 14658 5958 14660 6010
rect 14840 5958 14842 6010
rect 14596 5956 14602 5958
rect 14658 5956 14682 5958
rect 14738 5956 14762 5958
rect 14818 5956 14842 5958
rect 14898 5956 14904 5958
rect 14596 5936 14904 5956
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5370 11836 5510
rect 11867 5468 12175 5488
rect 11867 5466 11873 5468
rect 11929 5466 11953 5468
rect 12009 5466 12033 5468
rect 12089 5466 12113 5468
rect 12169 5466 12175 5468
rect 11929 5414 11931 5466
rect 12111 5414 12113 5466
rect 11867 5412 11873 5414
rect 11929 5412 11953 5414
rect 12009 5412 12033 5414
rect 12089 5412 12113 5414
rect 12169 5412 12175 5414
rect 11867 5392 12175 5412
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8772 2854 8800 2994
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 9138 2748 9446 2768
rect 9138 2746 9144 2748
rect 9200 2746 9224 2748
rect 9280 2746 9304 2748
rect 9360 2746 9384 2748
rect 9440 2746 9446 2748
rect 9200 2694 9202 2746
rect 9382 2694 9384 2746
rect 9138 2692 9144 2694
rect 9200 2692 9224 2694
rect 9280 2692 9304 2694
rect 9360 2692 9384 2694
rect 9440 2692 9446 2694
rect 9138 2672 9446 2692
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8220 2310 8248 2382
rect 9692 2378 9720 3606
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 3126 9812 3334
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10060 2514 10088 4014
rect 10980 4010 11008 5102
rect 11072 4146 11100 5170
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10244 3534 10272 3946
rect 11072 3738 11100 4082
rect 11808 4078 11836 5102
rect 13096 4622 13124 5646
rect 14596 4924 14904 4944
rect 14596 4922 14602 4924
rect 14658 4922 14682 4924
rect 14738 4922 14762 4924
rect 14818 4922 14842 4924
rect 14898 4922 14904 4924
rect 14658 4870 14660 4922
rect 14840 4870 14842 4922
rect 14596 4868 14602 4870
rect 14658 4868 14682 4870
rect 14738 4868 14762 4870
rect 14818 4868 14842 4870
rect 14898 4868 14904 4870
rect 14596 4848 14904 4868
rect 15764 4622 15792 17478
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 11867 4380 12175 4400
rect 11867 4378 11873 4380
rect 11929 4378 11953 4380
rect 12009 4378 12033 4380
rect 12089 4378 12113 4380
rect 12169 4378 12175 4380
rect 11929 4326 11931 4378
rect 12111 4326 12113 4378
rect 11867 4324 11873 4326
rect 11929 4324 11953 4326
rect 12009 4324 12033 4326
rect 12089 4324 12113 4326
rect 12169 4324 12175 4326
rect 11867 4304 12175 4324
rect 12912 4214 12940 4558
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14476 4214 14504 4422
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 2938 10272 3470
rect 11532 3466 11560 3878
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 10324 2984 10376 2990
rect 10244 2932 10324 2938
rect 10244 2926 10376 2932
rect 10244 2910 10364 2926
rect 10244 2650 10272 2910
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10796 2446 10824 2790
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 10428 800 10456 2314
rect 10796 2310 10824 2382
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 11808 2106 11836 4014
rect 12820 3738 12848 4014
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 11867 3292 12175 3312
rect 11867 3290 11873 3292
rect 11929 3290 11953 3292
rect 12009 3290 12033 3292
rect 12089 3290 12113 3292
rect 12169 3290 12175 3292
rect 11929 3238 11931 3290
rect 12111 3238 12113 3290
rect 11867 3236 11873 3238
rect 11929 3236 11953 3238
rect 12009 3236 12033 3238
rect 12089 3236 12113 3238
rect 12169 3236 12175 3238
rect 11867 3216 12175 3236
rect 12268 3074 12296 3674
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12176 3046 12296 3074
rect 12176 2514 12204 3046
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12268 2650 12296 2926
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12360 2582 12388 3538
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12452 2446 12480 3538
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 2650 12572 3334
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12544 2446 12572 2586
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 11867 2204 12175 2224
rect 11867 2202 11873 2204
rect 11929 2202 11953 2204
rect 12009 2202 12033 2204
rect 12089 2202 12113 2204
rect 12169 2202 12175 2204
rect 11929 2150 11931 2202
rect 12111 2150 12113 2202
rect 11867 2148 11873 2150
rect 11929 2148 11953 2150
rect 12009 2148 12033 2150
rect 12089 2148 12113 2150
rect 12169 2148 12175 2150
rect 11867 2128 12175 2148
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 12728 800 12756 3402
rect 12820 2446 12848 3470
rect 12912 3398 12940 4150
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14596 3836 14904 3856
rect 14596 3834 14602 3836
rect 14658 3834 14682 3836
rect 14738 3834 14762 3836
rect 14818 3834 14842 3836
rect 14898 3834 14904 3836
rect 14658 3782 14660 3834
rect 14840 3782 14842 3834
rect 14596 3780 14602 3782
rect 14658 3780 14682 3782
rect 14738 3780 14762 3782
rect 14818 3780 14842 3782
rect 14898 3780 14904 3782
rect 14596 3760 14904 3780
rect 14936 3534 14964 3878
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3126 12940 3334
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13096 2514 13124 3470
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 13360 2440 13412 2446
rect 13740 2394 13768 2790
rect 14292 2650 14320 3402
rect 14596 2748 14904 2768
rect 14596 2746 14602 2748
rect 14658 2746 14682 2748
rect 14738 2746 14762 2748
rect 14818 2746 14842 2748
rect 14898 2746 14904 2748
rect 14658 2694 14660 2746
rect 14840 2694 14842 2746
rect 14596 2692 14602 2694
rect 14658 2692 14682 2694
rect 14738 2692 14762 2694
rect 14818 2692 14842 2694
rect 14898 2692 14904 2694
rect 14596 2672 14904 2692
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14936 2446 14964 3470
rect 13412 2388 13768 2394
rect 13360 2382 13768 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 13372 2366 13768 2382
rect 13740 2310 13768 2366
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14108 2106 14136 2382
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 17316 2372 17368 2378
rect 17316 2314 17368 2320
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 15028 800 15056 2314
rect 17328 800 17356 2314
rect 1122 0 1178 800
rect 3422 0 3478 800
rect 5722 0 5778 800
rect 8022 0 8078 800
rect 10414 0 10470 800
rect 12714 0 12770 800
rect 15014 0 15070 800
rect 17314 0 17370 800
<< via2 >>
rect 6414 18522 6470 18524
rect 6494 18522 6550 18524
rect 6574 18522 6630 18524
rect 6654 18522 6710 18524
rect 6414 18470 6460 18522
rect 6460 18470 6470 18522
rect 6494 18470 6524 18522
rect 6524 18470 6536 18522
rect 6536 18470 6550 18522
rect 6574 18470 6588 18522
rect 6588 18470 6600 18522
rect 6600 18470 6630 18522
rect 6654 18470 6664 18522
rect 6664 18470 6710 18522
rect 6414 18468 6470 18470
rect 6494 18468 6550 18470
rect 6574 18468 6630 18470
rect 6654 18468 6710 18470
rect 3685 17978 3741 17980
rect 3765 17978 3821 17980
rect 3845 17978 3901 17980
rect 3925 17978 3981 17980
rect 3685 17926 3731 17978
rect 3731 17926 3741 17978
rect 3765 17926 3795 17978
rect 3795 17926 3807 17978
rect 3807 17926 3821 17978
rect 3845 17926 3859 17978
rect 3859 17926 3871 17978
rect 3871 17926 3901 17978
rect 3925 17926 3935 17978
rect 3935 17926 3981 17978
rect 3685 17924 3741 17926
rect 3765 17924 3821 17926
rect 3845 17924 3901 17926
rect 3925 17924 3981 17926
rect 11873 18522 11929 18524
rect 11953 18522 12009 18524
rect 12033 18522 12089 18524
rect 12113 18522 12169 18524
rect 11873 18470 11919 18522
rect 11919 18470 11929 18522
rect 11953 18470 11983 18522
rect 11983 18470 11995 18522
rect 11995 18470 12009 18522
rect 12033 18470 12047 18522
rect 12047 18470 12059 18522
rect 12059 18470 12089 18522
rect 12113 18470 12123 18522
rect 12123 18470 12169 18522
rect 11873 18468 11929 18470
rect 11953 18468 12009 18470
rect 12033 18468 12089 18470
rect 12113 18468 12169 18470
rect 9144 17978 9200 17980
rect 9224 17978 9280 17980
rect 9304 17978 9360 17980
rect 9384 17978 9440 17980
rect 9144 17926 9190 17978
rect 9190 17926 9200 17978
rect 9224 17926 9254 17978
rect 9254 17926 9266 17978
rect 9266 17926 9280 17978
rect 9304 17926 9318 17978
rect 9318 17926 9330 17978
rect 9330 17926 9360 17978
rect 9384 17926 9394 17978
rect 9394 17926 9440 17978
rect 9144 17924 9200 17926
rect 9224 17924 9280 17926
rect 9304 17924 9360 17926
rect 9384 17924 9440 17926
rect 6414 17434 6470 17436
rect 6494 17434 6550 17436
rect 6574 17434 6630 17436
rect 6654 17434 6710 17436
rect 6414 17382 6460 17434
rect 6460 17382 6470 17434
rect 6494 17382 6524 17434
rect 6524 17382 6536 17434
rect 6536 17382 6550 17434
rect 6574 17382 6588 17434
rect 6588 17382 6600 17434
rect 6600 17382 6630 17434
rect 6654 17382 6664 17434
rect 6664 17382 6710 17434
rect 6414 17380 6470 17382
rect 6494 17380 6550 17382
rect 6574 17380 6630 17382
rect 6654 17380 6710 17382
rect 3685 16890 3741 16892
rect 3765 16890 3821 16892
rect 3845 16890 3901 16892
rect 3925 16890 3981 16892
rect 3685 16838 3731 16890
rect 3731 16838 3741 16890
rect 3765 16838 3795 16890
rect 3795 16838 3807 16890
rect 3807 16838 3821 16890
rect 3845 16838 3859 16890
rect 3859 16838 3871 16890
rect 3871 16838 3901 16890
rect 3925 16838 3935 16890
rect 3935 16838 3981 16890
rect 3685 16836 3741 16838
rect 3765 16836 3821 16838
rect 3845 16836 3901 16838
rect 3925 16836 3981 16838
rect 9144 16890 9200 16892
rect 9224 16890 9280 16892
rect 9304 16890 9360 16892
rect 9384 16890 9440 16892
rect 9144 16838 9190 16890
rect 9190 16838 9200 16890
rect 9224 16838 9254 16890
rect 9254 16838 9266 16890
rect 9266 16838 9280 16890
rect 9304 16838 9318 16890
rect 9318 16838 9330 16890
rect 9330 16838 9360 16890
rect 9384 16838 9394 16890
rect 9394 16838 9440 16890
rect 9144 16836 9200 16838
rect 9224 16836 9280 16838
rect 9304 16836 9360 16838
rect 9384 16836 9440 16838
rect 6414 16346 6470 16348
rect 6494 16346 6550 16348
rect 6574 16346 6630 16348
rect 6654 16346 6710 16348
rect 6414 16294 6460 16346
rect 6460 16294 6470 16346
rect 6494 16294 6524 16346
rect 6524 16294 6536 16346
rect 6536 16294 6550 16346
rect 6574 16294 6588 16346
rect 6588 16294 6600 16346
rect 6600 16294 6630 16346
rect 6654 16294 6664 16346
rect 6664 16294 6710 16346
rect 6414 16292 6470 16294
rect 6494 16292 6550 16294
rect 6574 16292 6630 16294
rect 6654 16292 6710 16294
rect 3685 15802 3741 15804
rect 3765 15802 3821 15804
rect 3845 15802 3901 15804
rect 3925 15802 3981 15804
rect 3685 15750 3731 15802
rect 3731 15750 3741 15802
rect 3765 15750 3795 15802
rect 3795 15750 3807 15802
rect 3807 15750 3821 15802
rect 3845 15750 3859 15802
rect 3859 15750 3871 15802
rect 3871 15750 3901 15802
rect 3925 15750 3935 15802
rect 3935 15750 3981 15802
rect 3685 15748 3741 15750
rect 3765 15748 3821 15750
rect 3845 15748 3901 15750
rect 3925 15748 3981 15750
rect 9144 15802 9200 15804
rect 9224 15802 9280 15804
rect 9304 15802 9360 15804
rect 9384 15802 9440 15804
rect 9144 15750 9190 15802
rect 9190 15750 9200 15802
rect 9224 15750 9254 15802
rect 9254 15750 9266 15802
rect 9266 15750 9280 15802
rect 9304 15750 9318 15802
rect 9318 15750 9330 15802
rect 9330 15750 9360 15802
rect 9384 15750 9394 15802
rect 9394 15750 9440 15802
rect 9144 15748 9200 15750
rect 9224 15748 9280 15750
rect 9304 15748 9360 15750
rect 9384 15748 9440 15750
rect 6414 15258 6470 15260
rect 6494 15258 6550 15260
rect 6574 15258 6630 15260
rect 6654 15258 6710 15260
rect 6414 15206 6460 15258
rect 6460 15206 6470 15258
rect 6494 15206 6524 15258
rect 6524 15206 6536 15258
rect 6536 15206 6550 15258
rect 6574 15206 6588 15258
rect 6588 15206 6600 15258
rect 6600 15206 6630 15258
rect 6654 15206 6664 15258
rect 6664 15206 6710 15258
rect 6414 15204 6470 15206
rect 6494 15204 6550 15206
rect 6574 15204 6630 15206
rect 6654 15204 6710 15206
rect 3685 14714 3741 14716
rect 3765 14714 3821 14716
rect 3845 14714 3901 14716
rect 3925 14714 3981 14716
rect 3685 14662 3731 14714
rect 3731 14662 3741 14714
rect 3765 14662 3795 14714
rect 3795 14662 3807 14714
rect 3807 14662 3821 14714
rect 3845 14662 3859 14714
rect 3859 14662 3871 14714
rect 3871 14662 3901 14714
rect 3925 14662 3935 14714
rect 3935 14662 3981 14714
rect 3685 14660 3741 14662
rect 3765 14660 3821 14662
rect 3845 14660 3901 14662
rect 3925 14660 3981 14662
rect 9144 14714 9200 14716
rect 9224 14714 9280 14716
rect 9304 14714 9360 14716
rect 9384 14714 9440 14716
rect 9144 14662 9190 14714
rect 9190 14662 9200 14714
rect 9224 14662 9254 14714
rect 9254 14662 9266 14714
rect 9266 14662 9280 14714
rect 9304 14662 9318 14714
rect 9318 14662 9330 14714
rect 9330 14662 9360 14714
rect 9384 14662 9394 14714
rect 9394 14662 9440 14714
rect 9144 14660 9200 14662
rect 9224 14660 9280 14662
rect 9304 14660 9360 14662
rect 9384 14660 9440 14662
rect 6414 14170 6470 14172
rect 6494 14170 6550 14172
rect 6574 14170 6630 14172
rect 6654 14170 6710 14172
rect 6414 14118 6460 14170
rect 6460 14118 6470 14170
rect 6494 14118 6524 14170
rect 6524 14118 6536 14170
rect 6536 14118 6550 14170
rect 6574 14118 6588 14170
rect 6588 14118 6600 14170
rect 6600 14118 6630 14170
rect 6654 14118 6664 14170
rect 6664 14118 6710 14170
rect 6414 14116 6470 14118
rect 6494 14116 6550 14118
rect 6574 14116 6630 14118
rect 6654 14116 6710 14118
rect 3685 13626 3741 13628
rect 3765 13626 3821 13628
rect 3845 13626 3901 13628
rect 3925 13626 3981 13628
rect 3685 13574 3731 13626
rect 3731 13574 3741 13626
rect 3765 13574 3795 13626
rect 3795 13574 3807 13626
rect 3807 13574 3821 13626
rect 3845 13574 3859 13626
rect 3859 13574 3871 13626
rect 3871 13574 3901 13626
rect 3925 13574 3935 13626
rect 3935 13574 3981 13626
rect 3685 13572 3741 13574
rect 3765 13572 3821 13574
rect 3845 13572 3901 13574
rect 3925 13572 3981 13574
rect 9144 13626 9200 13628
rect 9224 13626 9280 13628
rect 9304 13626 9360 13628
rect 9384 13626 9440 13628
rect 9144 13574 9190 13626
rect 9190 13574 9200 13626
rect 9224 13574 9254 13626
rect 9254 13574 9266 13626
rect 9266 13574 9280 13626
rect 9304 13574 9318 13626
rect 9318 13574 9330 13626
rect 9330 13574 9360 13626
rect 9384 13574 9394 13626
rect 9394 13574 9440 13626
rect 9144 13572 9200 13574
rect 9224 13572 9280 13574
rect 9304 13572 9360 13574
rect 9384 13572 9440 13574
rect 6414 13082 6470 13084
rect 6494 13082 6550 13084
rect 6574 13082 6630 13084
rect 6654 13082 6710 13084
rect 6414 13030 6460 13082
rect 6460 13030 6470 13082
rect 6494 13030 6524 13082
rect 6524 13030 6536 13082
rect 6536 13030 6550 13082
rect 6574 13030 6588 13082
rect 6588 13030 6600 13082
rect 6600 13030 6630 13082
rect 6654 13030 6664 13082
rect 6664 13030 6710 13082
rect 6414 13028 6470 13030
rect 6494 13028 6550 13030
rect 6574 13028 6630 13030
rect 6654 13028 6710 13030
rect 3685 12538 3741 12540
rect 3765 12538 3821 12540
rect 3845 12538 3901 12540
rect 3925 12538 3981 12540
rect 3685 12486 3731 12538
rect 3731 12486 3741 12538
rect 3765 12486 3795 12538
rect 3795 12486 3807 12538
rect 3807 12486 3821 12538
rect 3845 12486 3859 12538
rect 3859 12486 3871 12538
rect 3871 12486 3901 12538
rect 3925 12486 3935 12538
rect 3935 12486 3981 12538
rect 3685 12484 3741 12486
rect 3765 12484 3821 12486
rect 3845 12484 3901 12486
rect 3925 12484 3981 12486
rect 9144 12538 9200 12540
rect 9224 12538 9280 12540
rect 9304 12538 9360 12540
rect 9384 12538 9440 12540
rect 9144 12486 9190 12538
rect 9190 12486 9200 12538
rect 9224 12486 9254 12538
rect 9254 12486 9266 12538
rect 9266 12486 9280 12538
rect 9304 12486 9318 12538
rect 9318 12486 9330 12538
rect 9330 12486 9360 12538
rect 9384 12486 9394 12538
rect 9394 12486 9440 12538
rect 9144 12484 9200 12486
rect 9224 12484 9280 12486
rect 9304 12484 9360 12486
rect 9384 12484 9440 12486
rect 6414 11994 6470 11996
rect 6494 11994 6550 11996
rect 6574 11994 6630 11996
rect 6654 11994 6710 11996
rect 6414 11942 6460 11994
rect 6460 11942 6470 11994
rect 6494 11942 6524 11994
rect 6524 11942 6536 11994
rect 6536 11942 6550 11994
rect 6574 11942 6588 11994
rect 6588 11942 6600 11994
rect 6600 11942 6630 11994
rect 6654 11942 6664 11994
rect 6664 11942 6710 11994
rect 6414 11940 6470 11942
rect 6494 11940 6550 11942
rect 6574 11940 6630 11942
rect 6654 11940 6710 11942
rect 3685 11450 3741 11452
rect 3765 11450 3821 11452
rect 3845 11450 3901 11452
rect 3925 11450 3981 11452
rect 3685 11398 3731 11450
rect 3731 11398 3741 11450
rect 3765 11398 3795 11450
rect 3795 11398 3807 11450
rect 3807 11398 3821 11450
rect 3845 11398 3859 11450
rect 3859 11398 3871 11450
rect 3871 11398 3901 11450
rect 3925 11398 3935 11450
rect 3935 11398 3981 11450
rect 3685 11396 3741 11398
rect 3765 11396 3821 11398
rect 3845 11396 3901 11398
rect 3925 11396 3981 11398
rect 9144 11450 9200 11452
rect 9224 11450 9280 11452
rect 9304 11450 9360 11452
rect 9384 11450 9440 11452
rect 9144 11398 9190 11450
rect 9190 11398 9200 11450
rect 9224 11398 9254 11450
rect 9254 11398 9266 11450
rect 9266 11398 9280 11450
rect 9304 11398 9318 11450
rect 9318 11398 9330 11450
rect 9330 11398 9360 11450
rect 9384 11398 9394 11450
rect 9394 11398 9440 11450
rect 9144 11396 9200 11398
rect 9224 11396 9280 11398
rect 9304 11396 9360 11398
rect 9384 11396 9440 11398
rect 6414 10906 6470 10908
rect 6494 10906 6550 10908
rect 6574 10906 6630 10908
rect 6654 10906 6710 10908
rect 6414 10854 6460 10906
rect 6460 10854 6470 10906
rect 6494 10854 6524 10906
rect 6524 10854 6536 10906
rect 6536 10854 6550 10906
rect 6574 10854 6588 10906
rect 6588 10854 6600 10906
rect 6600 10854 6630 10906
rect 6654 10854 6664 10906
rect 6664 10854 6710 10906
rect 6414 10852 6470 10854
rect 6494 10852 6550 10854
rect 6574 10852 6630 10854
rect 6654 10852 6710 10854
rect 3685 10362 3741 10364
rect 3765 10362 3821 10364
rect 3845 10362 3901 10364
rect 3925 10362 3981 10364
rect 3685 10310 3731 10362
rect 3731 10310 3741 10362
rect 3765 10310 3795 10362
rect 3795 10310 3807 10362
rect 3807 10310 3821 10362
rect 3845 10310 3859 10362
rect 3859 10310 3871 10362
rect 3871 10310 3901 10362
rect 3925 10310 3935 10362
rect 3935 10310 3981 10362
rect 3685 10308 3741 10310
rect 3765 10308 3821 10310
rect 3845 10308 3901 10310
rect 3925 10308 3981 10310
rect 9144 10362 9200 10364
rect 9224 10362 9280 10364
rect 9304 10362 9360 10364
rect 9384 10362 9440 10364
rect 9144 10310 9190 10362
rect 9190 10310 9200 10362
rect 9224 10310 9254 10362
rect 9254 10310 9266 10362
rect 9266 10310 9280 10362
rect 9304 10310 9318 10362
rect 9318 10310 9330 10362
rect 9330 10310 9360 10362
rect 9384 10310 9394 10362
rect 9394 10310 9440 10362
rect 9144 10308 9200 10310
rect 9224 10308 9280 10310
rect 9304 10308 9360 10310
rect 9384 10308 9440 10310
rect 6414 9818 6470 9820
rect 6494 9818 6550 9820
rect 6574 9818 6630 9820
rect 6654 9818 6710 9820
rect 6414 9766 6460 9818
rect 6460 9766 6470 9818
rect 6494 9766 6524 9818
rect 6524 9766 6536 9818
rect 6536 9766 6550 9818
rect 6574 9766 6588 9818
rect 6588 9766 6600 9818
rect 6600 9766 6630 9818
rect 6654 9766 6664 9818
rect 6664 9766 6710 9818
rect 6414 9764 6470 9766
rect 6494 9764 6550 9766
rect 6574 9764 6630 9766
rect 6654 9764 6710 9766
rect 3685 9274 3741 9276
rect 3765 9274 3821 9276
rect 3845 9274 3901 9276
rect 3925 9274 3981 9276
rect 3685 9222 3731 9274
rect 3731 9222 3741 9274
rect 3765 9222 3795 9274
rect 3795 9222 3807 9274
rect 3807 9222 3821 9274
rect 3845 9222 3859 9274
rect 3859 9222 3871 9274
rect 3871 9222 3901 9274
rect 3925 9222 3935 9274
rect 3935 9222 3981 9274
rect 3685 9220 3741 9222
rect 3765 9220 3821 9222
rect 3845 9220 3901 9222
rect 3925 9220 3981 9222
rect 9144 9274 9200 9276
rect 9224 9274 9280 9276
rect 9304 9274 9360 9276
rect 9384 9274 9440 9276
rect 9144 9222 9190 9274
rect 9190 9222 9200 9274
rect 9224 9222 9254 9274
rect 9254 9222 9266 9274
rect 9266 9222 9280 9274
rect 9304 9222 9318 9274
rect 9318 9222 9330 9274
rect 9330 9222 9360 9274
rect 9384 9222 9394 9274
rect 9394 9222 9440 9274
rect 9144 9220 9200 9222
rect 9224 9220 9280 9222
rect 9304 9220 9360 9222
rect 9384 9220 9440 9222
rect 6414 8730 6470 8732
rect 6494 8730 6550 8732
rect 6574 8730 6630 8732
rect 6654 8730 6710 8732
rect 6414 8678 6460 8730
rect 6460 8678 6470 8730
rect 6494 8678 6524 8730
rect 6524 8678 6536 8730
rect 6536 8678 6550 8730
rect 6574 8678 6588 8730
rect 6588 8678 6600 8730
rect 6600 8678 6630 8730
rect 6654 8678 6664 8730
rect 6664 8678 6710 8730
rect 6414 8676 6470 8678
rect 6494 8676 6550 8678
rect 6574 8676 6630 8678
rect 6654 8676 6710 8678
rect 3685 8186 3741 8188
rect 3765 8186 3821 8188
rect 3845 8186 3901 8188
rect 3925 8186 3981 8188
rect 3685 8134 3731 8186
rect 3731 8134 3741 8186
rect 3765 8134 3795 8186
rect 3795 8134 3807 8186
rect 3807 8134 3821 8186
rect 3845 8134 3859 8186
rect 3859 8134 3871 8186
rect 3871 8134 3901 8186
rect 3925 8134 3935 8186
rect 3935 8134 3981 8186
rect 3685 8132 3741 8134
rect 3765 8132 3821 8134
rect 3845 8132 3901 8134
rect 3925 8132 3981 8134
rect 9144 8186 9200 8188
rect 9224 8186 9280 8188
rect 9304 8186 9360 8188
rect 9384 8186 9440 8188
rect 9144 8134 9190 8186
rect 9190 8134 9200 8186
rect 9224 8134 9254 8186
rect 9254 8134 9266 8186
rect 9266 8134 9280 8186
rect 9304 8134 9318 8186
rect 9318 8134 9330 8186
rect 9330 8134 9360 8186
rect 9384 8134 9394 8186
rect 9394 8134 9440 8186
rect 9144 8132 9200 8134
rect 9224 8132 9280 8134
rect 9304 8132 9360 8134
rect 9384 8132 9440 8134
rect 6414 7642 6470 7644
rect 6494 7642 6550 7644
rect 6574 7642 6630 7644
rect 6654 7642 6710 7644
rect 6414 7590 6460 7642
rect 6460 7590 6470 7642
rect 6494 7590 6524 7642
rect 6524 7590 6536 7642
rect 6536 7590 6550 7642
rect 6574 7590 6588 7642
rect 6588 7590 6600 7642
rect 6600 7590 6630 7642
rect 6654 7590 6664 7642
rect 6664 7590 6710 7642
rect 6414 7588 6470 7590
rect 6494 7588 6550 7590
rect 6574 7588 6630 7590
rect 6654 7588 6710 7590
rect 3685 7098 3741 7100
rect 3765 7098 3821 7100
rect 3845 7098 3901 7100
rect 3925 7098 3981 7100
rect 3685 7046 3731 7098
rect 3731 7046 3741 7098
rect 3765 7046 3795 7098
rect 3795 7046 3807 7098
rect 3807 7046 3821 7098
rect 3845 7046 3859 7098
rect 3859 7046 3871 7098
rect 3871 7046 3901 7098
rect 3925 7046 3935 7098
rect 3935 7046 3981 7098
rect 3685 7044 3741 7046
rect 3765 7044 3821 7046
rect 3845 7044 3901 7046
rect 3925 7044 3981 7046
rect 9144 7098 9200 7100
rect 9224 7098 9280 7100
rect 9304 7098 9360 7100
rect 9384 7098 9440 7100
rect 9144 7046 9190 7098
rect 9190 7046 9200 7098
rect 9224 7046 9254 7098
rect 9254 7046 9266 7098
rect 9266 7046 9280 7098
rect 9304 7046 9318 7098
rect 9318 7046 9330 7098
rect 9330 7046 9360 7098
rect 9384 7046 9394 7098
rect 9394 7046 9440 7098
rect 9144 7044 9200 7046
rect 9224 7044 9280 7046
rect 9304 7044 9360 7046
rect 9384 7044 9440 7046
rect 6414 6554 6470 6556
rect 6494 6554 6550 6556
rect 6574 6554 6630 6556
rect 6654 6554 6710 6556
rect 6414 6502 6460 6554
rect 6460 6502 6470 6554
rect 6494 6502 6524 6554
rect 6524 6502 6536 6554
rect 6536 6502 6550 6554
rect 6574 6502 6588 6554
rect 6588 6502 6600 6554
rect 6600 6502 6630 6554
rect 6654 6502 6664 6554
rect 6664 6502 6710 6554
rect 6414 6500 6470 6502
rect 6494 6500 6550 6502
rect 6574 6500 6630 6502
rect 6654 6500 6710 6502
rect 3685 6010 3741 6012
rect 3765 6010 3821 6012
rect 3845 6010 3901 6012
rect 3925 6010 3981 6012
rect 3685 5958 3731 6010
rect 3731 5958 3741 6010
rect 3765 5958 3795 6010
rect 3795 5958 3807 6010
rect 3807 5958 3821 6010
rect 3845 5958 3859 6010
rect 3859 5958 3871 6010
rect 3871 5958 3901 6010
rect 3925 5958 3935 6010
rect 3935 5958 3981 6010
rect 3685 5956 3741 5958
rect 3765 5956 3821 5958
rect 3845 5956 3901 5958
rect 3925 5956 3981 5958
rect 9144 6010 9200 6012
rect 9224 6010 9280 6012
rect 9304 6010 9360 6012
rect 9384 6010 9440 6012
rect 9144 5958 9190 6010
rect 9190 5958 9200 6010
rect 9224 5958 9254 6010
rect 9254 5958 9266 6010
rect 9266 5958 9280 6010
rect 9304 5958 9318 6010
rect 9318 5958 9330 6010
rect 9330 5958 9360 6010
rect 9384 5958 9394 6010
rect 9394 5958 9440 6010
rect 9144 5956 9200 5958
rect 9224 5956 9280 5958
rect 9304 5956 9360 5958
rect 9384 5956 9440 5958
rect 6414 5466 6470 5468
rect 6494 5466 6550 5468
rect 6574 5466 6630 5468
rect 6654 5466 6710 5468
rect 6414 5414 6460 5466
rect 6460 5414 6470 5466
rect 6494 5414 6524 5466
rect 6524 5414 6536 5466
rect 6536 5414 6550 5466
rect 6574 5414 6588 5466
rect 6588 5414 6600 5466
rect 6600 5414 6630 5466
rect 6654 5414 6664 5466
rect 6664 5414 6710 5466
rect 6414 5412 6470 5414
rect 6494 5412 6550 5414
rect 6574 5412 6630 5414
rect 6654 5412 6710 5414
rect 3685 4922 3741 4924
rect 3765 4922 3821 4924
rect 3845 4922 3901 4924
rect 3925 4922 3981 4924
rect 3685 4870 3731 4922
rect 3731 4870 3741 4922
rect 3765 4870 3795 4922
rect 3795 4870 3807 4922
rect 3807 4870 3821 4922
rect 3845 4870 3859 4922
rect 3859 4870 3871 4922
rect 3871 4870 3901 4922
rect 3925 4870 3935 4922
rect 3935 4870 3981 4922
rect 3685 4868 3741 4870
rect 3765 4868 3821 4870
rect 3845 4868 3901 4870
rect 3925 4868 3981 4870
rect 6414 4378 6470 4380
rect 6494 4378 6550 4380
rect 6574 4378 6630 4380
rect 6654 4378 6710 4380
rect 6414 4326 6460 4378
rect 6460 4326 6470 4378
rect 6494 4326 6524 4378
rect 6524 4326 6536 4378
rect 6536 4326 6550 4378
rect 6574 4326 6588 4378
rect 6588 4326 6600 4378
rect 6600 4326 6630 4378
rect 6654 4326 6664 4378
rect 6664 4326 6710 4378
rect 6414 4324 6470 4326
rect 6494 4324 6550 4326
rect 6574 4324 6630 4326
rect 6654 4324 6710 4326
rect 3685 3834 3741 3836
rect 3765 3834 3821 3836
rect 3845 3834 3901 3836
rect 3925 3834 3981 3836
rect 3685 3782 3731 3834
rect 3731 3782 3741 3834
rect 3765 3782 3795 3834
rect 3795 3782 3807 3834
rect 3807 3782 3821 3834
rect 3845 3782 3859 3834
rect 3859 3782 3871 3834
rect 3871 3782 3901 3834
rect 3925 3782 3935 3834
rect 3935 3782 3981 3834
rect 3685 3780 3741 3782
rect 3765 3780 3821 3782
rect 3845 3780 3901 3782
rect 3925 3780 3981 3782
rect 6414 3290 6470 3292
rect 6494 3290 6550 3292
rect 6574 3290 6630 3292
rect 6654 3290 6710 3292
rect 6414 3238 6460 3290
rect 6460 3238 6470 3290
rect 6494 3238 6524 3290
rect 6524 3238 6536 3290
rect 6536 3238 6550 3290
rect 6574 3238 6588 3290
rect 6588 3238 6600 3290
rect 6600 3238 6630 3290
rect 6654 3238 6664 3290
rect 6664 3238 6710 3290
rect 6414 3236 6470 3238
rect 6494 3236 6550 3238
rect 6574 3236 6630 3238
rect 6654 3236 6710 3238
rect 3685 2746 3741 2748
rect 3765 2746 3821 2748
rect 3845 2746 3901 2748
rect 3925 2746 3981 2748
rect 3685 2694 3731 2746
rect 3731 2694 3741 2746
rect 3765 2694 3795 2746
rect 3795 2694 3807 2746
rect 3807 2694 3821 2746
rect 3845 2694 3859 2746
rect 3859 2694 3871 2746
rect 3871 2694 3901 2746
rect 3925 2694 3935 2746
rect 3935 2694 3981 2746
rect 3685 2692 3741 2694
rect 3765 2692 3821 2694
rect 3845 2692 3901 2694
rect 3925 2692 3981 2694
rect 6414 2202 6470 2204
rect 6494 2202 6550 2204
rect 6574 2202 6630 2204
rect 6654 2202 6710 2204
rect 6414 2150 6460 2202
rect 6460 2150 6470 2202
rect 6494 2150 6524 2202
rect 6524 2150 6536 2202
rect 6536 2150 6550 2202
rect 6574 2150 6588 2202
rect 6588 2150 6600 2202
rect 6600 2150 6630 2202
rect 6654 2150 6664 2202
rect 6664 2150 6710 2202
rect 6414 2148 6470 2150
rect 6494 2148 6550 2150
rect 6574 2148 6630 2150
rect 6654 2148 6710 2150
rect 9144 4922 9200 4924
rect 9224 4922 9280 4924
rect 9304 4922 9360 4924
rect 9384 4922 9440 4924
rect 9144 4870 9190 4922
rect 9190 4870 9200 4922
rect 9224 4870 9254 4922
rect 9254 4870 9266 4922
rect 9266 4870 9280 4922
rect 9304 4870 9318 4922
rect 9318 4870 9330 4922
rect 9330 4870 9360 4922
rect 9384 4870 9394 4922
rect 9394 4870 9440 4922
rect 9144 4868 9200 4870
rect 9224 4868 9280 4870
rect 9304 4868 9360 4870
rect 9384 4868 9440 4870
rect 9144 3834 9200 3836
rect 9224 3834 9280 3836
rect 9304 3834 9360 3836
rect 9384 3834 9440 3836
rect 9144 3782 9190 3834
rect 9190 3782 9200 3834
rect 9224 3782 9254 3834
rect 9254 3782 9266 3834
rect 9266 3782 9280 3834
rect 9304 3782 9318 3834
rect 9318 3782 9330 3834
rect 9330 3782 9360 3834
rect 9384 3782 9394 3834
rect 9394 3782 9440 3834
rect 9144 3780 9200 3782
rect 9224 3780 9280 3782
rect 9304 3780 9360 3782
rect 9384 3780 9440 3782
rect 14602 17978 14658 17980
rect 14682 17978 14738 17980
rect 14762 17978 14818 17980
rect 14842 17978 14898 17980
rect 14602 17926 14648 17978
rect 14648 17926 14658 17978
rect 14682 17926 14712 17978
rect 14712 17926 14724 17978
rect 14724 17926 14738 17978
rect 14762 17926 14776 17978
rect 14776 17926 14788 17978
rect 14788 17926 14818 17978
rect 14842 17926 14852 17978
rect 14852 17926 14898 17978
rect 14602 17924 14658 17926
rect 14682 17924 14738 17926
rect 14762 17924 14818 17926
rect 14842 17924 14898 17926
rect 11873 17434 11929 17436
rect 11953 17434 12009 17436
rect 12033 17434 12089 17436
rect 12113 17434 12169 17436
rect 11873 17382 11919 17434
rect 11919 17382 11929 17434
rect 11953 17382 11983 17434
rect 11983 17382 11995 17434
rect 11995 17382 12009 17434
rect 12033 17382 12047 17434
rect 12047 17382 12059 17434
rect 12059 17382 12089 17434
rect 12113 17382 12123 17434
rect 12123 17382 12169 17434
rect 11873 17380 11929 17382
rect 11953 17380 12009 17382
rect 12033 17380 12089 17382
rect 12113 17380 12169 17382
rect 14602 16890 14658 16892
rect 14682 16890 14738 16892
rect 14762 16890 14818 16892
rect 14842 16890 14898 16892
rect 14602 16838 14648 16890
rect 14648 16838 14658 16890
rect 14682 16838 14712 16890
rect 14712 16838 14724 16890
rect 14724 16838 14738 16890
rect 14762 16838 14776 16890
rect 14776 16838 14788 16890
rect 14788 16838 14818 16890
rect 14842 16838 14852 16890
rect 14852 16838 14898 16890
rect 14602 16836 14658 16838
rect 14682 16836 14738 16838
rect 14762 16836 14818 16838
rect 14842 16836 14898 16838
rect 11873 16346 11929 16348
rect 11953 16346 12009 16348
rect 12033 16346 12089 16348
rect 12113 16346 12169 16348
rect 11873 16294 11919 16346
rect 11919 16294 11929 16346
rect 11953 16294 11983 16346
rect 11983 16294 11995 16346
rect 11995 16294 12009 16346
rect 12033 16294 12047 16346
rect 12047 16294 12059 16346
rect 12059 16294 12089 16346
rect 12113 16294 12123 16346
rect 12123 16294 12169 16346
rect 11873 16292 11929 16294
rect 11953 16292 12009 16294
rect 12033 16292 12089 16294
rect 12113 16292 12169 16294
rect 14602 15802 14658 15804
rect 14682 15802 14738 15804
rect 14762 15802 14818 15804
rect 14842 15802 14898 15804
rect 14602 15750 14648 15802
rect 14648 15750 14658 15802
rect 14682 15750 14712 15802
rect 14712 15750 14724 15802
rect 14724 15750 14738 15802
rect 14762 15750 14776 15802
rect 14776 15750 14788 15802
rect 14788 15750 14818 15802
rect 14842 15750 14852 15802
rect 14852 15750 14898 15802
rect 14602 15748 14658 15750
rect 14682 15748 14738 15750
rect 14762 15748 14818 15750
rect 14842 15748 14898 15750
rect 11873 15258 11929 15260
rect 11953 15258 12009 15260
rect 12033 15258 12089 15260
rect 12113 15258 12169 15260
rect 11873 15206 11919 15258
rect 11919 15206 11929 15258
rect 11953 15206 11983 15258
rect 11983 15206 11995 15258
rect 11995 15206 12009 15258
rect 12033 15206 12047 15258
rect 12047 15206 12059 15258
rect 12059 15206 12089 15258
rect 12113 15206 12123 15258
rect 12123 15206 12169 15258
rect 11873 15204 11929 15206
rect 11953 15204 12009 15206
rect 12033 15204 12089 15206
rect 12113 15204 12169 15206
rect 14602 14714 14658 14716
rect 14682 14714 14738 14716
rect 14762 14714 14818 14716
rect 14842 14714 14898 14716
rect 14602 14662 14648 14714
rect 14648 14662 14658 14714
rect 14682 14662 14712 14714
rect 14712 14662 14724 14714
rect 14724 14662 14738 14714
rect 14762 14662 14776 14714
rect 14776 14662 14788 14714
rect 14788 14662 14818 14714
rect 14842 14662 14852 14714
rect 14852 14662 14898 14714
rect 14602 14660 14658 14662
rect 14682 14660 14738 14662
rect 14762 14660 14818 14662
rect 14842 14660 14898 14662
rect 11873 14170 11929 14172
rect 11953 14170 12009 14172
rect 12033 14170 12089 14172
rect 12113 14170 12169 14172
rect 11873 14118 11919 14170
rect 11919 14118 11929 14170
rect 11953 14118 11983 14170
rect 11983 14118 11995 14170
rect 11995 14118 12009 14170
rect 12033 14118 12047 14170
rect 12047 14118 12059 14170
rect 12059 14118 12089 14170
rect 12113 14118 12123 14170
rect 12123 14118 12169 14170
rect 11873 14116 11929 14118
rect 11953 14116 12009 14118
rect 12033 14116 12089 14118
rect 12113 14116 12169 14118
rect 14602 13626 14658 13628
rect 14682 13626 14738 13628
rect 14762 13626 14818 13628
rect 14842 13626 14898 13628
rect 14602 13574 14648 13626
rect 14648 13574 14658 13626
rect 14682 13574 14712 13626
rect 14712 13574 14724 13626
rect 14724 13574 14738 13626
rect 14762 13574 14776 13626
rect 14776 13574 14788 13626
rect 14788 13574 14818 13626
rect 14842 13574 14852 13626
rect 14852 13574 14898 13626
rect 14602 13572 14658 13574
rect 14682 13572 14738 13574
rect 14762 13572 14818 13574
rect 14842 13572 14898 13574
rect 11873 13082 11929 13084
rect 11953 13082 12009 13084
rect 12033 13082 12089 13084
rect 12113 13082 12169 13084
rect 11873 13030 11919 13082
rect 11919 13030 11929 13082
rect 11953 13030 11983 13082
rect 11983 13030 11995 13082
rect 11995 13030 12009 13082
rect 12033 13030 12047 13082
rect 12047 13030 12059 13082
rect 12059 13030 12089 13082
rect 12113 13030 12123 13082
rect 12123 13030 12169 13082
rect 11873 13028 11929 13030
rect 11953 13028 12009 13030
rect 12033 13028 12089 13030
rect 12113 13028 12169 13030
rect 14602 12538 14658 12540
rect 14682 12538 14738 12540
rect 14762 12538 14818 12540
rect 14842 12538 14898 12540
rect 14602 12486 14648 12538
rect 14648 12486 14658 12538
rect 14682 12486 14712 12538
rect 14712 12486 14724 12538
rect 14724 12486 14738 12538
rect 14762 12486 14776 12538
rect 14776 12486 14788 12538
rect 14788 12486 14818 12538
rect 14842 12486 14852 12538
rect 14852 12486 14898 12538
rect 14602 12484 14658 12486
rect 14682 12484 14738 12486
rect 14762 12484 14818 12486
rect 14842 12484 14898 12486
rect 11873 11994 11929 11996
rect 11953 11994 12009 11996
rect 12033 11994 12089 11996
rect 12113 11994 12169 11996
rect 11873 11942 11919 11994
rect 11919 11942 11929 11994
rect 11953 11942 11983 11994
rect 11983 11942 11995 11994
rect 11995 11942 12009 11994
rect 12033 11942 12047 11994
rect 12047 11942 12059 11994
rect 12059 11942 12089 11994
rect 12113 11942 12123 11994
rect 12123 11942 12169 11994
rect 11873 11940 11929 11942
rect 11953 11940 12009 11942
rect 12033 11940 12089 11942
rect 12113 11940 12169 11942
rect 14602 11450 14658 11452
rect 14682 11450 14738 11452
rect 14762 11450 14818 11452
rect 14842 11450 14898 11452
rect 14602 11398 14648 11450
rect 14648 11398 14658 11450
rect 14682 11398 14712 11450
rect 14712 11398 14724 11450
rect 14724 11398 14738 11450
rect 14762 11398 14776 11450
rect 14776 11398 14788 11450
rect 14788 11398 14818 11450
rect 14842 11398 14852 11450
rect 14852 11398 14898 11450
rect 14602 11396 14658 11398
rect 14682 11396 14738 11398
rect 14762 11396 14818 11398
rect 14842 11396 14898 11398
rect 11873 10906 11929 10908
rect 11953 10906 12009 10908
rect 12033 10906 12089 10908
rect 12113 10906 12169 10908
rect 11873 10854 11919 10906
rect 11919 10854 11929 10906
rect 11953 10854 11983 10906
rect 11983 10854 11995 10906
rect 11995 10854 12009 10906
rect 12033 10854 12047 10906
rect 12047 10854 12059 10906
rect 12059 10854 12089 10906
rect 12113 10854 12123 10906
rect 12123 10854 12169 10906
rect 11873 10852 11929 10854
rect 11953 10852 12009 10854
rect 12033 10852 12089 10854
rect 12113 10852 12169 10854
rect 14602 10362 14658 10364
rect 14682 10362 14738 10364
rect 14762 10362 14818 10364
rect 14842 10362 14898 10364
rect 14602 10310 14648 10362
rect 14648 10310 14658 10362
rect 14682 10310 14712 10362
rect 14712 10310 14724 10362
rect 14724 10310 14738 10362
rect 14762 10310 14776 10362
rect 14776 10310 14788 10362
rect 14788 10310 14818 10362
rect 14842 10310 14852 10362
rect 14852 10310 14898 10362
rect 14602 10308 14658 10310
rect 14682 10308 14738 10310
rect 14762 10308 14818 10310
rect 14842 10308 14898 10310
rect 11873 9818 11929 9820
rect 11953 9818 12009 9820
rect 12033 9818 12089 9820
rect 12113 9818 12169 9820
rect 11873 9766 11919 9818
rect 11919 9766 11929 9818
rect 11953 9766 11983 9818
rect 11983 9766 11995 9818
rect 11995 9766 12009 9818
rect 12033 9766 12047 9818
rect 12047 9766 12059 9818
rect 12059 9766 12089 9818
rect 12113 9766 12123 9818
rect 12123 9766 12169 9818
rect 11873 9764 11929 9766
rect 11953 9764 12009 9766
rect 12033 9764 12089 9766
rect 12113 9764 12169 9766
rect 14602 9274 14658 9276
rect 14682 9274 14738 9276
rect 14762 9274 14818 9276
rect 14842 9274 14898 9276
rect 14602 9222 14648 9274
rect 14648 9222 14658 9274
rect 14682 9222 14712 9274
rect 14712 9222 14724 9274
rect 14724 9222 14738 9274
rect 14762 9222 14776 9274
rect 14776 9222 14788 9274
rect 14788 9222 14818 9274
rect 14842 9222 14852 9274
rect 14852 9222 14898 9274
rect 14602 9220 14658 9222
rect 14682 9220 14738 9222
rect 14762 9220 14818 9222
rect 14842 9220 14898 9222
rect 11873 8730 11929 8732
rect 11953 8730 12009 8732
rect 12033 8730 12089 8732
rect 12113 8730 12169 8732
rect 11873 8678 11919 8730
rect 11919 8678 11929 8730
rect 11953 8678 11983 8730
rect 11983 8678 11995 8730
rect 11995 8678 12009 8730
rect 12033 8678 12047 8730
rect 12047 8678 12059 8730
rect 12059 8678 12089 8730
rect 12113 8678 12123 8730
rect 12123 8678 12169 8730
rect 11873 8676 11929 8678
rect 11953 8676 12009 8678
rect 12033 8676 12089 8678
rect 12113 8676 12169 8678
rect 14602 8186 14658 8188
rect 14682 8186 14738 8188
rect 14762 8186 14818 8188
rect 14842 8186 14898 8188
rect 14602 8134 14648 8186
rect 14648 8134 14658 8186
rect 14682 8134 14712 8186
rect 14712 8134 14724 8186
rect 14724 8134 14738 8186
rect 14762 8134 14776 8186
rect 14776 8134 14788 8186
rect 14788 8134 14818 8186
rect 14842 8134 14852 8186
rect 14852 8134 14898 8186
rect 14602 8132 14658 8134
rect 14682 8132 14738 8134
rect 14762 8132 14818 8134
rect 14842 8132 14898 8134
rect 11873 7642 11929 7644
rect 11953 7642 12009 7644
rect 12033 7642 12089 7644
rect 12113 7642 12169 7644
rect 11873 7590 11919 7642
rect 11919 7590 11929 7642
rect 11953 7590 11983 7642
rect 11983 7590 11995 7642
rect 11995 7590 12009 7642
rect 12033 7590 12047 7642
rect 12047 7590 12059 7642
rect 12059 7590 12089 7642
rect 12113 7590 12123 7642
rect 12123 7590 12169 7642
rect 11873 7588 11929 7590
rect 11953 7588 12009 7590
rect 12033 7588 12089 7590
rect 12113 7588 12169 7590
rect 14602 7098 14658 7100
rect 14682 7098 14738 7100
rect 14762 7098 14818 7100
rect 14842 7098 14898 7100
rect 14602 7046 14648 7098
rect 14648 7046 14658 7098
rect 14682 7046 14712 7098
rect 14712 7046 14724 7098
rect 14724 7046 14738 7098
rect 14762 7046 14776 7098
rect 14776 7046 14788 7098
rect 14788 7046 14818 7098
rect 14842 7046 14852 7098
rect 14852 7046 14898 7098
rect 14602 7044 14658 7046
rect 14682 7044 14738 7046
rect 14762 7044 14818 7046
rect 14842 7044 14898 7046
rect 11873 6554 11929 6556
rect 11953 6554 12009 6556
rect 12033 6554 12089 6556
rect 12113 6554 12169 6556
rect 11873 6502 11919 6554
rect 11919 6502 11929 6554
rect 11953 6502 11983 6554
rect 11983 6502 11995 6554
rect 11995 6502 12009 6554
rect 12033 6502 12047 6554
rect 12047 6502 12059 6554
rect 12059 6502 12089 6554
rect 12113 6502 12123 6554
rect 12123 6502 12169 6554
rect 11873 6500 11929 6502
rect 11953 6500 12009 6502
rect 12033 6500 12089 6502
rect 12113 6500 12169 6502
rect 14602 6010 14658 6012
rect 14682 6010 14738 6012
rect 14762 6010 14818 6012
rect 14842 6010 14898 6012
rect 14602 5958 14648 6010
rect 14648 5958 14658 6010
rect 14682 5958 14712 6010
rect 14712 5958 14724 6010
rect 14724 5958 14738 6010
rect 14762 5958 14776 6010
rect 14776 5958 14788 6010
rect 14788 5958 14818 6010
rect 14842 5958 14852 6010
rect 14852 5958 14898 6010
rect 14602 5956 14658 5958
rect 14682 5956 14738 5958
rect 14762 5956 14818 5958
rect 14842 5956 14898 5958
rect 11873 5466 11929 5468
rect 11953 5466 12009 5468
rect 12033 5466 12089 5468
rect 12113 5466 12169 5468
rect 11873 5414 11919 5466
rect 11919 5414 11929 5466
rect 11953 5414 11983 5466
rect 11983 5414 11995 5466
rect 11995 5414 12009 5466
rect 12033 5414 12047 5466
rect 12047 5414 12059 5466
rect 12059 5414 12089 5466
rect 12113 5414 12123 5466
rect 12123 5414 12169 5466
rect 11873 5412 11929 5414
rect 11953 5412 12009 5414
rect 12033 5412 12089 5414
rect 12113 5412 12169 5414
rect 9144 2746 9200 2748
rect 9224 2746 9280 2748
rect 9304 2746 9360 2748
rect 9384 2746 9440 2748
rect 9144 2694 9190 2746
rect 9190 2694 9200 2746
rect 9224 2694 9254 2746
rect 9254 2694 9266 2746
rect 9266 2694 9280 2746
rect 9304 2694 9318 2746
rect 9318 2694 9330 2746
rect 9330 2694 9360 2746
rect 9384 2694 9394 2746
rect 9394 2694 9440 2746
rect 9144 2692 9200 2694
rect 9224 2692 9280 2694
rect 9304 2692 9360 2694
rect 9384 2692 9440 2694
rect 14602 4922 14658 4924
rect 14682 4922 14738 4924
rect 14762 4922 14818 4924
rect 14842 4922 14898 4924
rect 14602 4870 14648 4922
rect 14648 4870 14658 4922
rect 14682 4870 14712 4922
rect 14712 4870 14724 4922
rect 14724 4870 14738 4922
rect 14762 4870 14776 4922
rect 14776 4870 14788 4922
rect 14788 4870 14818 4922
rect 14842 4870 14852 4922
rect 14852 4870 14898 4922
rect 14602 4868 14658 4870
rect 14682 4868 14738 4870
rect 14762 4868 14818 4870
rect 14842 4868 14898 4870
rect 11873 4378 11929 4380
rect 11953 4378 12009 4380
rect 12033 4378 12089 4380
rect 12113 4378 12169 4380
rect 11873 4326 11919 4378
rect 11919 4326 11929 4378
rect 11953 4326 11983 4378
rect 11983 4326 11995 4378
rect 11995 4326 12009 4378
rect 12033 4326 12047 4378
rect 12047 4326 12059 4378
rect 12059 4326 12089 4378
rect 12113 4326 12123 4378
rect 12123 4326 12169 4378
rect 11873 4324 11929 4326
rect 11953 4324 12009 4326
rect 12033 4324 12089 4326
rect 12113 4324 12169 4326
rect 11873 3290 11929 3292
rect 11953 3290 12009 3292
rect 12033 3290 12089 3292
rect 12113 3290 12169 3292
rect 11873 3238 11919 3290
rect 11919 3238 11929 3290
rect 11953 3238 11983 3290
rect 11983 3238 11995 3290
rect 11995 3238 12009 3290
rect 12033 3238 12047 3290
rect 12047 3238 12059 3290
rect 12059 3238 12089 3290
rect 12113 3238 12123 3290
rect 12123 3238 12169 3290
rect 11873 3236 11929 3238
rect 11953 3236 12009 3238
rect 12033 3236 12089 3238
rect 12113 3236 12169 3238
rect 11873 2202 11929 2204
rect 11953 2202 12009 2204
rect 12033 2202 12089 2204
rect 12113 2202 12169 2204
rect 11873 2150 11919 2202
rect 11919 2150 11929 2202
rect 11953 2150 11983 2202
rect 11983 2150 11995 2202
rect 11995 2150 12009 2202
rect 12033 2150 12047 2202
rect 12047 2150 12059 2202
rect 12059 2150 12089 2202
rect 12113 2150 12123 2202
rect 12123 2150 12169 2202
rect 11873 2148 11929 2150
rect 11953 2148 12009 2150
rect 12033 2148 12089 2150
rect 12113 2148 12169 2150
rect 14602 3834 14658 3836
rect 14682 3834 14738 3836
rect 14762 3834 14818 3836
rect 14842 3834 14898 3836
rect 14602 3782 14648 3834
rect 14648 3782 14658 3834
rect 14682 3782 14712 3834
rect 14712 3782 14724 3834
rect 14724 3782 14738 3834
rect 14762 3782 14776 3834
rect 14776 3782 14788 3834
rect 14788 3782 14818 3834
rect 14842 3782 14852 3834
rect 14852 3782 14898 3834
rect 14602 3780 14658 3782
rect 14682 3780 14738 3782
rect 14762 3780 14818 3782
rect 14842 3780 14898 3782
rect 14602 2746 14658 2748
rect 14682 2746 14738 2748
rect 14762 2746 14818 2748
rect 14842 2746 14898 2748
rect 14602 2694 14648 2746
rect 14648 2694 14658 2746
rect 14682 2694 14712 2746
rect 14712 2694 14724 2746
rect 14724 2694 14738 2746
rect 14762 2694 14776 2746
rect 14776 2694 14788 2746
rect 14788 2694 14818 2746
rect 14842 2694 14852 2746
rect 14852 2694 14898 2746
rect 14602 2692 14658 2694
rect 14682 2692 14738 2694
rect 14762 2692 14818 2694
rect 14842 2692 14898 2694
<< metal3 >>
rect 6402 18528 6722 18529
rect 6402 18464 6410 18528
rect 6474 18464 6490 18528
rect 6554 18464 6570 18528
rect 6634 18464 6650 18528
rect 6714 18464 6722 18528
rect 6402 18463 6722 18464
rect 11861 18528 12181 18529
rect 11861 18464 11869 18528
rect 11933 18464 11949 18528
rect 12013 18464 12029 18528
rect 12093 18464 12109 18528
rect 12173 18464 12181 18528
rect 11861 18463 12181 18464
rect 3673 17984 3993 17985
rect 3673 17920 3681 17984
rect 3745 17920 3761 17984
rect 3825 17920 3841 17984
rect 3905 17920 3921 17984
rect 3985 17920 3993 17984
rect 3673 17919 3993 17920
rect 9132 17984 9452 17985
rect 9132 17920 9140 17984
rect 9204 17920 9220 17984
rect 9284 17920 9300 17984
rect 9364 17920 9380 17984
rect 9444 17920 9452 17984
rect 9132 17919 9452 17920
rect 14590 17984 14910 17985
rect 14590 17920 14598 17984
rect 14662 17920 14678 17984
rect 14742 17920 14758 17984
rect 14822 17920 14838 17984
rect 14902 17920 14910 17984
rect 14590 17919 14910 17920
rect 6402 17440 6722 17441
rect 6402 17376 6410 17440
rect 6474 17376 6490 17440
rect 6554 17376 6570 17440
rect 6634 17376 6650 17440
rect 6714 17376 6722 17440
rect 6402 17375 6722 17376
rect 11861 17440 12181 17441
rect 11861 17376 11869 17440
rect 11933 17376 11949 17440
rect 12013 17376 12029 17440
rect 12093 17376 12109 17440
rect 12173 17376 12181 17440
rect 11861 17375 12181 17376
rect 3673 16896 3993 16897
rect 3673 16832 3681 16896
rect 3745 16832 3761 16896
rect 3825 16832 3841 16896
rect 3905 16832 3921 16896
rect 3985 16832 3993 16896
rect 3673 16831 3993 16832
rect 9132 16896 9452 16897
rect 9132 16832 9140 16896
rect 9204 16832 9220 16896
rect 9284 16832 9300 16896
rect 9364 16832 9380 16896
rect 9444 16832 9452 16896
rect 9132 16831 9452 16832
rect 14590 16896 14910 16897
rect 14590 16832 14598 16896
rect 14662 16832 14678 16896
rect 14742 16832 14758 16896
rect 14822 16832 14838 16896
rect 14902 16832 14910 16896
rect 14590 16831 14910 16832
rect 6402 16352 6722 16353
rect 6402 16288 6410 16352
rect 6474 16288 6490 16352
rect 6554 16288 6570 16352
rect 6634 16288 6650 16352
rect 6714 16288 6722 16352
rect 6402 16287 6722 16288
rect 11861 16352 12181 16353
rect 11861 16288 11869 16352
rect 11933 16288 11949 16352
rect 12013 16288 12029 16352
rect 12093 16288 12109 16352
rect 12173 16288 12181 16352
rect 11861 16287 12181 16288
rect 3673 15808 3993 15809
rect 3673 15744 3681 15808
rect 3745 15744 3761 15808
rect 3825 15744 3841 15808
rect 3905 15744 3921 15808
rect 3985 15744 3993 15808
rect 3673 15743 3993 15744
rect 9132 15808 9452 15809
rect 9132 15744 9140 15808
rect 9204 15744 9220 15808
rect 9284 15744 9300 15808
rect 9364 15744 9380 15808
rect 9444 15744 9452 15808
rect 9132 15743 9452 15744
rect 14590 15808 14910 15809
rect 14590 15744 14598 15808
rect 14662 15744 14678 15808
rect 14742 15744 14758 15808
rect 14822 15744 14838 15808
rect 14902 15744 14910 15808
rect 14590 15743 14910 15744
rect 6402 15264 6722 15265
rect 6402 15200 6410 15264
rect 6474 15200 6490 15264
rect 6554 15200 6570 15264
rect 6634 15200 6650 15264
rect 6714 15200 6722 15264
rect 6402 15199 6722 15200
rect 11861 15264 12181 15265
rect 11861 15200 11869 15264
rect 11933 15200 11949 15264
rect 12013 15200 12029 15264
rect 12093 15200 12109 15264
rect 12173 15200 12181 15264
rect 11861 15199 12181 15200
rect 3673 14720 3993 14721
rect 3673 14656 3681 14720
rect 3745 14656 3761 14720
rect 3825 14656 3841 14720
rect 3905 14656 3921 14720
rect 3985 14656 3993 14720
rect 3673 14655 3993 14656
rect 9132 14720 9452 14721
rect 9132 14656 9140 14720
rect 9204 14656 9220 14720
rect 9284 14656 9300 14720
rect 9364 14656 9380 14720
rect 9444 14656 9452 14720
rect 9132 14655 9452 14656
rect 14590 14720 14910 14721
rect 14590 14656 14598 14720
rect 14662 14656 14678 14720
rect 14742 14656 14758 14720
rect 14822 14656 14838 14720
rect 14902 14656 14910 14720
rect 14590 14655 14910 14656
rect 6402 14176 6722 14177
rect 6402 14112 6410 14176
rect 6474 14112 6490 14176
rect 6554 14112 6570 14176
rect 6634 14112 6650 14176
rect 6714 14112 6722 14176
rect 6402 14111 6722 14112
rect 11861 14176 12181 14177
rect 11861 14112 11869 14176
rect 11933 14112 11949 14176
rect 12013 14112 12029 14176
rect 12093 14112 12109 14176
rect 12173 14112 12181 14176
rect 11861 14111 12181 14112
rect 3673 13632 3993 13633
rect 3673 13568 3681 13632
rect 3745 13568 3761 13632
rect 3825 13568 3841 13632
rect 3905 13568 3921 13632
rect 3985 13568 3993 13632
rect 3673 13567 3993 13568
rect 9132 13632 9452 13633
rect 9132 13568 9140 13632
rect 9204 13568 9220 13632
rect 9284 13568 9300 13632
rect 9364 13568 9380 13632
rect 9444 13568 9452 13632
rect 9132 13567 9452 13568
rect 14590 13632 14910 13633
rect 14590 13568 14598 13632
rect 14662 13568 14678 13632
rect 14742 13568 14758 13632
rect 14822 13568 14838 13632
rect 14902 13568 14910 13632
rect 14590 13567 14910 13568
rect 6402 13088 6722 13089
rect 6402 13024 6410 13088
rect 6474 13024 6490 13088
rect 6554 13024 6570 13088
rect 6634 13024 6650 13088
rect 6714 13024 6722 13088
rect 6402 13023 6722 13024
rect 11861 13088 12181 13089
rect 11861 13024 11869 13088
rect 11933 13024 11949 13088
rect 12013 13024 12029 13088
rect 12093 13024 12109 13088
rect 12173 13024 12181 13088
rect 11861 13023 12181 13024
rect 3673 12544 3993 12545
rect 3673 12480 3681 12544
rect 3745 12480 3761 12544
rect 3825 12480 3841 12544
rect 3905 12480 3921 12544
rect 3985 12480 3993 12544
rect 3673 12479 3993 12480
rect 9132 12544 9452 12545
rect 9132 12480 9140 12544
rect 9204 12480 9220 12544
rect 9284 12480 9300 12544
rect 9364 12480 9380 12544
rect 9444 12480 9452 12544
rect 9132 12479 9452 12480
rect 14590 12544 14910 12545
rect 14590 12480 14598 12544
rect 14662 12480 14678 12544
rect 14742 12480 14758 12544
rect 14822 12480 14838 12544
rect 14902 12480 14910 12544
rect 14590 12479 14910 12480
rect 6402 12000 6722 12001
rect 6402 11936 6410 12000
rect 6474 11936 6490 12000
rect 6554 11936 6570 12000
rect 6634 11936 6650 12000
rect 6714 11936 6722 12000
rect 6402 11935 6722 11936
rect 11861 12000 12181 12001
rect 11861 11936 11869 12000
rect 11933 11936 11949 12000
rect 12013 11936 12029 12000
rect 12093 11936 12109 12000
rect 12173 11936 12181 12000
rect 11861 11935 12181 11936
rect 3673 11456 3993 11457
rect 3673 11392 3681 11456
rect 3745 11392 3761 11456
rect 3825 11392 3841 11456
rect 3905 11392 3921 11456
rect 3985 11392 3993 11456
rect 3673 11391 3993 11392
rect 9132 11456 9452 11457
rect 9132 11392 9140 11456
rect 9204 11392 9220 11456
rect 9284 11392 9300 11456
rect 9364 11392 9380 11456
rect 9444 11392 9452 11456
rect 9132 11391 9452 11392
rect 14590 11456 14910 11457
rect 14590 11392 14598 11456
rect 14662 11392 14678 11456
rect 14742 11392 14758 11456
rect 14822 11392 14838 11456
rect 14902 11392 14910 11456
rect 14590 11391 14910 11392
rect 6402 10912 6722 10913
rect 6402 10848 6410 10912
rect 6474 10848 6490 10912
rect 6554 10848 6570 10912
rect 6634 10848 6650 10912
rect 6714 10848 6722 10912
rect 6402 10847 6722 10848
rect 11861 10912 12181 10913
rect 11861 10848 11869 10912
rect 11933 10848 11949 10912
rect 12013 10848 12029 10912
rect 12093 10848 12109 10912
rect 12173 10848 12181 10912
rect 11861 10847 12181 10848
rect 3673 10368 3993 10369
rect 3673 10304 3681 10368
rect 3745 10304 3761 10368
rect 3825 10304 3841 10368
rect 3905 10304 3921 10368
rect 3985 10304 3993 10368
rect 3673 10303 3993 10304
rect 9132 10368 9452 10369
rect 9132 10304 9140 10368
rect 9204 10304 9220 10368
rect 9284 10304 9300 10368
rect 9364 10304 9380 10368
rect 9444 10304 9452 10368
rect 9132 10303 9452 10304
rect 14590 10368 14910 10369
rect 14590 10304 14598 10368
rect 14662 10304 14678 10368
rect 14742 10304 14758 10368
rect 14822 10304 14838 10368
rect 14902 10304 14910 10368
rect 14590 10303 14910 10304
rect 6402 9824 6722 9825
rect 6402 9760 6410 9824
rect 6474 9760 6490 9824
rect 6554 9760 6570 9824
rect 6634 9760 6650 9824
rect 6714 9760 6722 9824
rect 6402 9759 6722 9760
rect 11861 9824 12181 9825
rect 11861 9760 11869 9824
rect 11933 9760 11949 9824
rect 12013 9760 12029 9824
rect 12093 9760 12109 9824
rect 12173 9760 12181 9824
rect 11861 9759 12181 9760
rect 3673 9280 3993 9281
rect 3673 9216 3681 9280
rect 3745 9216 3761 9280
rect 3825 9216 3841 9280
rect 3905 9216 3921 9280
rect 3985 9216 3993 9280
rect 3673 9215 3993 9216
rect 9132 9280 9452 9281
rect 9132 9216 9140 9280
rect 9204 9216 9220 9280
rect 9284 9216 9300 9280
rect 9364 9216 9380 9280
rect 9444 9216 9452 9280
rect 9132 9215 9452 9216
rect 14590 9280 14910 9281
rect 14590 9216 14598 9280
rect 14662 9216 14678 9280
rect 14742 9216 14758 9280
rect 14822 9216 14838 9280
rect 14902 9216 14910 9280
rect 14590 9215 14910 9216
rect 6402 8736 6722 8737
rect 6402 8672 6410 8736
rect 6474 8672 6490 8736
rect 6554 8672 6570 8736
rect 6634 8672 6650 8736
rect 6714 8672 6722 8736
rect 6402 8671 6722 8672
rect 11861 8736 12181 8737
rect 11861 8672 11869 8736
rect 11933 8672 11949 8736
rect 12013 8672 12029 8736
rect 12093 8672 12109 8736
rect 12173 8672 12181 8736
rect 11861 8671 12181 8672
rect 3673 8192 3993 8193
rect 3673 8128 3681 8192
rect 3745 8128 3761 8192
rect 3825 8128 3841 8192
rect 3905 8128 3921 8192
rect 3985 8128 3993 8192
rect 3673 8127 3993 8128
rect 9132 8192 9452 8193
rect 9132 8128 9140 8192
rect 9204 8128 9220 8192
rect 9284 8128 9300 8192
rect 9364 8128 9380 8192
rect 9444 8128 9452 8192
rect 9132 8127 9452 8128
rect 14590 8192 14910 8193
rect 14590 8128 14598 8192
rect 14662 8128 14678 8192
rect 14742 8128 14758 8192
rect 14822 8128 14838 8192
rect 14902 8128 14910 8192
rect 14590 8127 14910 8128
rect 6402 7648 6722 7649
rect 6402 7584 6410 7648
rect 6474 7584 6490 7648
rect 6554 7584 6570 7648
rect 6634 7584 6650 7648
rect 6714 7584 6722 7648
rect 6402 7583 6722 7584
rect 11861 7648 12181 7649
rect 11861 7584 11869 7648
rect 11933 7584 11949 7648
rect 12013 7584 12029 7648
rect 12093 7584 12109 7648
rect 12173 7584 12181 7648
rect 11861 7583 12181 7584
rect 3673 7104 3993 7105
rect 3673 7040 3681 7104
rect 3745 7040 3761 7104
rect 3825 7040 3841 7104
rect 3905 7040 3921 7104
rect 3985 7040 3993 7104
rect 3673 7039 3993 7040
rect 9132 7104 9452 7105
rect 9132 7040 9140 7104
rect 9204 7040 9220 7104
rect 9284 7040 9300 7104
rect 9364 7040 9380 7104
rect 9444 7040 9452 7104
rect 9132 7039 9452 7040
rect 14590 7104 14910 7105
rect 14590 7040 14598 7104
rect 14662 7040 14678 7104
rect 14742 7040 14758 7104
rect 14822 7040 14838 7104
rect 14902 7040 14910 7104
rect 14590 7039 14910 7040
rect 6402 6560 6722 6561
rect 6402 6496 6410 6560
rect 6474 6496 6490 6560
rect 6554 6496 6570 6560
rect 6634 6496 6650 6560
rect 6714 6496 6722 6560
rect 6402 6495 6722 6496
rect 11861 6560 12181 6561
rect 11861 6496 11869 6560
rect 11933 6496 11949 6560
rect 12013 6496 12029 6560
rect 12093 6496 12109 6560
rect 12173 6496 12181 6560
rect 11861 6495 12181 6496
rect 3673 6016 3993 6017
rect 3673 5952 3681 6016
rect 3745 5952 3761 6016
rect 3825 5952 3841 6016
rect 3905 5952 3921 6016
rect 3985 5952 3993 6016
rect 3673 5951 3993 5952
rect 9132 6016 9452 6017
rect 9132 5952 9140 6016
rect 9204 5952 9220 6016
rect 9284 5952 9300 6016
rect 9364 5952 9380 6016
rect 9444 5952 9452 6016
rect 9132 5951 9452 5952
rect 14590 6016 14910 6017
rect 14590 5952 14598 6016
rect 14662 5952 14678 6016
rect 14742 5952 14758 6016
rect 14822 5952 14838 6016
rect 14902 5952 14910 6016
rect 14590 5951 14910 5952
rect 6402 5472 6722 5473
rect 6402 5408 6410 5472
rect 6474 5408 6490 5472
rect 6554 5408 6570 5472
rect 6634 5408 6650 5472
rect 6714 5408 6722 5472
rect 6402 5407 6722 5408
rect 11861 5472 12181 5473
rect 11861 5408 11869 5472
rect 11933 5408 11949 5472
rect 12013 5408 12029 5472
rect 12093 5408 12109 5472
rect 12173 5408 12181 5472
rect 11861 5407 12181 5408
rect 3673 4928 3993 4929
rect 3673 4864 3681 4928
rect 3745 4864 3761 4928
rect 3825 4864 3841 4928
rect 3905 4864 3921 4928
rect 3985 4864 3993 4928
rect 3673 4863 3993 4864
rect 9132 4928 9452 4929
rect 9132 4864 9140 4928
rect 9204 4864 9220 4928
rect 9284 4864 9300 4928
rect 9364 4864 9380 4928
rect 9444 4864 9452 4928
rect 9132 4863 9452 4864
rect 14590 4928 14910 4929
rect 14590 4864 14598 4928
rect 14662 4864 14678 4928
rect 14742 4864 14758 4928
rect 14822 4864 14838 4928
rect 14902 4864 14910 4928
rect 14590 4863 14910 4864
rect 6402 4384 6722 4385
rect 6402 4320 6410 4384
rect 6474 4320 6490 4384
rect 6554 4320 6570 4384
rect 6634 4320 6650 4384
rect 6714 4320 6722 4384
rect 6402 4319 6722 4320
rect 11861 4384 12181 4385
rect 11861 4320 11869 4384
rect 11933 4320 11949 4384
rect 12013 4320 12029 4384
rect 12093 4320 12109 4384
rect 12173 4320 12181 4384
rect 11861 4319 12181 4320
rect 3673 3840 3993 3841
rect 3673 3776 3681 3840
rect 3745 3776 3761 3840
rect 3825 3776 3841 3840
rect 3905 3776 3921 3840
rect 3985 3776 3993 3840
rect 3673 3775 3993 3776
rect 9132 3840 9452 3841
rect 9132 3776 9140 3840
rect 9204 3776 9220 3840
rect 9284 3776 9300 3840
rect 9364 3776 9380 3840
rect 9444 3776 9452 3840
rect 9132 3775 9452 3776
rect 14590 3840 14910 3841
rect 14590 3776 14598 3840
rect 14662 3776 14678 3840
rect 14742 3776 14758 3840
rect 14822 3776 14838 3840
rect 14902 3776 14910 3840
rect 14590 3775 14910 3776
rect 6402 3296 6722 3297
rect 6402 3232 6410 3296
rect 6474 3232 6490 3296
rect 6554 3232 6570 3296
rect 6634 3232 6650 3296
rect 6714 3232 6722 3296
rect 6402 3231 6722 3232
rect 11861 3296 12181 3297
rect 11861 3232 11869 3296
rect 11933 3232 11949 3296
rect 12013 3232 12029 3296
rect 12093 3232 12109 3296
rect 12173 3232 12181 3296
rect 11861 3231 12181 3232
rect 3673 2752 3993 2753
rect 3673 2688 3681 2752
rect 3745 2688 3761 2752
rect 3825 2688 3841 2752
rect 3905 2688 3921 2752
rect 3985 2688 3993 2752
rect 3673 2687 3993 2688
rect 9132 2752 9452 2753
rect 9132 2688 9140 2752
rect 9204 2688 9220 2752
rect 9284 2688 9300 2752
rect 9364 2688 9380 2752
rect 9444 2688 9452 2752
rect 9132 2687 9452 2688
rect 14590 2752 14910 2753
rect 14590 2688 14598 2752
rect 14662 2688 14678 2752
rect 14742 2688 14758 2752
rect 14822 2688 14838 2752
rect 14902 2688 14910 2752
rect 14590 2687 14910 2688
rect 6402 2208 6722 2209
rect 6402 2144 6410 2208
rect 6474 2144 6490 2208
rect 6554 2144 6570 2208
rect 6634 2144 6650 2208
rect 6714 2144 6722 2208
rect 6402 2143 6722 2144
rect 11861 2208 12181 2209
rect 11861 2144 11869 2208
rect 11933 2144 11949 2208
rect 12013 2144 12029 2208
rect 12093 2144 12109 2208
rect 12173 2144 12181 2208
rect 11861 2143 12181 2144
<< via3 >>
rect 6410 18524 6474 18528
rect 6410 18468 6414 18524
rect 6414 18468 6470 18524
rect 6470 18468 6474 18524
rect 6410 18464 6474 18468
rect 6490 18524 6554 18528
rect 6490 18468 6494 18524
rect 6494 18468 6550 18524
rect 6550 18468 6554 18524
rect 6490 18464 6554 18468
rect 6570 18524 6634 18528
rect 6570 18468 6574 18524
rect 6574 18468 6630 18524
rect 6630 18468 6634 18524
rect 6570 18464 6634 18468
rect 6650 18524 6714 18528
rect 6650 18468 6654 18524
rect 6654 18468 6710 18524
rect 6710 18468 6714 18524
rect 6650 18464 6714 18468
rect 11869 18524 11933 18528
rect 11869 18468 11873 18524
rect 11873 18468 11929 18524
rect 11929 18468 11933 18524
rect 11869 18464 11933 18468
rect 11949 18524 12013 18528
rect 11949 18468 11953 18524
rect 11953 18468 12009 18524
rect 12009 18468 12013 18524
rect 11949 18464 12013 18468
rect 12029 18524 12093 18528
rect 12029 18468 12033 18524
rect 12033 18468 12089 18524
rect 12089 18468 12093 18524
rect 12029 18464 12093 18468
rect 12109 18524 12173 18528
rect 12109 18468 12113 18524
rect 12113 18468 12169 18524
rect 12169 18468 12173 18524
rect 12109 18464 12173 18468
rect 3681 17980 3745 17984
rect 3681 17924 3685 17980
rect 3685 17924 3741 17980
rect 3741 17924 3745 17980
rect 3681 17920 3745 17924
rect 3761 17980 3825 17984
rect 3761 17924 3765 17980
rect 3765 17924 3821 17980
rect 3821 17924 3825 17980
rect 3761 17920 3825 17924
rect 3841 17980 3905 17984
rect 3841 17924 3845 17980
rect 3845 17924 3901 17980
rect 3901 17924 3905 17980
rect 3841 17920 3905 17924
rect 3921 17980 3985 17984
rect 3921 17924 3925 17980
rect 3925 17924 3981 17980
rect 3981 17924 3985 17980
rect 3921 17920 3985 17924
rect 9140 17980 9204 17984
rect 9140 17924 9144 17980
rect 9144 17924 9200 17980
rect 9200 17924 9204 17980
rect 9140 17920 9204 17924
rect 9220 17980 9284 17984
rect 9220 17924 9224 17980
rect 9224 17924 9280 17980
rect 9280 17924 9284 17980
rect 9220 17920 9284 17924
rect 9300 17980 9364 17984
rect 9300 17924 9304 17980
rect 9304 17924 9360 17980
rect 9360 17924 9364 17980
rect 9300 17920 9364 17924
rect 9380 17980 9444 17984
rect 9380 17924 9384 17980
rect 9384 17924 9440 17980
rect 9440 17924 9444 17980
rect 9380 17920 9444 17924
rect 14598 17980 14662 17984
rect 14598 17924 14602 17980
rect 14602 17924 14658 17980
rect 14658 17924 14662 17980
rect 14598 17920 14662 17924
rect 14678 17980 14742 17984
rect 14678 17924 14682 17980
rect 14682 17924 14738 17980
rect 14738 17924 14742 17980
rect 14678 17920 14742 17924
rect 14758 17980 14822 17984
rect 14758 17924 14762 17980
rect 14762 17924 14818 17980
rect 14818 17924 14822 17980
rect 14758 17920 14822 17924
rect 14838 17980 14902 17984
rect 14838 17924 14842 17980
rect 14842 17924 14898 17980
rect 14898 17924 14902 17980
rect 14838 17920 14902 17924
rect 6410 17436 6474 17440
rect 6410 17380 6414 17436
rect 6414 17380 6470 17436
rect 6470 17380 6474 17436
rect 6410 17376 6474 17380
rect 6490 17436 6554 17440
rect 6490 17380 6494 17436
rect 6494 17380 6550 17436
rect 6550 17380 6554 17436
rect 6490 17376 6554 17380
rect 6570 17436 6634 17440
rect 6570 17380 6574 17436
rect 6574 17380 6630 17436
rect 6630 17380 6634 17436
rect 6570 17376 6634 17380
rect 6650 17436 6714 17440
rect 6650 17380 6654 17436
rect 6654 17380 6710 17436
rect 6710 17380 6714 17436
rect 6650 17376 6714 17380
rect 11869 17436 11933 17440
rect 11869 17380 11873 17436
rect 11873 17380 11929 17436
rect 11929 17380 11933 17436
rect 11869 17376 11933 17380
rect 11949 17436 12013 17440
rect 11949 17380 11953 17436
rect 11953 17380 12009 17436
rect 12009 17380 12013 17436
rect 11949 17376 12013 17380
rect 12029 17436 12093 17440
rect 12029 17380 12033 17436
rect 12033 17380 12089 17436
rect 12089 17380 12093 17436
rect 12029 17376 12093 17380
rect 12109 17436 12173 17440
rect 12109 17380 12113 17436
rect 12113 17380 12169 17436
rect 12169 17380 12173 17436
rect 12109 17376 12173 17380
rect 3681 16892 3745 16896
rect 3681 16836 3685 16892
rect 3685 16836 3741 16892
rect 3741 16836 3745 16892
rect 3681 16832 3745 16836
rect 3761 16892 3825 16896
rect 3761 16836 3765 16892
rect 3765 16836 3821 16892
rect 3821 16836 3825 16892
rect 3761 16832 3825 16836
rect 3841 16892 3905 16896
rect 3841 16836 3845 16892
rect 3845 16836 3901 16892
rect 3901 16836 3905 16892
rect 3841 16832 3905 16836
rect 3921 16892 3985 16896
rect 3921 16836 3925 16892
rect 3925 16836 3981 16892
rect 3981 16836 3985 16892
rect 3921 16832 3985 16836
rect 9140 16892 9204 16896
rect 9140 16836 9144 16892
rect 9144 16836 9200 16892
rect 9200 16836 9204 16892
rect 9140 16832 9204 16836
rect 9220 16892 9284 16896
rect 9220 16836 9224 16892
rect 9224 16836 9280 16892
rect 9280 16836 9284 16892
rect 9220 16832 9284 16836
rect 9300 16892 9364 16896
rect 9300 16836 9304 16892
rect 9304 16836 9360 16892
rect 9360 16836 9364 16892
rect 9300 16832 9364 16836
rect 9380 16892 9444 16896
rect 9380 16836 9384 16892
rect 9384 16836 9440 16892
rect 9440 16836 9444 16892
rect 9380 16832 9444 16836
rect 14598 16892 14662 16896
rect 14598 16836 14602 16892
rect 14602 16836 14658 16892
rect 14658 16836 14662 16892
rect 14598 16832 14662 16836
rect 14678 16892 14742 16896
rect 14678 16836 14682 16892
rect 14682 16836 14738 16892
rect 14738 16836 14742 16892
rect 14678 16832 14742 16836
rect 14758 16892 14822 16896
rect 14758 16836 14762 16892
rect 14762 16836 14818 16892
rect 14818 16836 14822 16892
rect 14758 16832 14822 16836
rect 14838 16892 14902 16896
rect 14838 16836 14842 16892
rect 14842 16836 14898 16892
rect 14898 16836 14902 16892
rect 14838 16832 14902 16836
rect 6410 16348 6474 16352
rect 6410 16292 6414 16348
rect 6414 16292 6470 16348
rect 6470 16292 6474 16348
rect 6410 16288 6474 16292
rect 6490 16348 6554 16352
rect 6490 16292 6494 16348
rect 6494 16292 6550 16348
rect 6550 16292 6554 16348
rect 6490 16288 6554 16292
rect 6570 16348 6634 16352
rect 6570 16292 6574 16348
rect 6574 16292 6630 16348
rect 6630 16292 6634 16348
rect 6570 16288 6634 16292
rect 6650 16348 6714 16352
rect 6650 16292 6654 16348
rect 6654 16292 6710 16348
rect 6710 16292 6714 16348
rect 6650 16288 6714 16292
rect 11869 16348 11933 16352
rect 11869 16292 11873 16348
rect 11873 16292 11929 16348
rect 11929 16292 11933 16348
rect 11869 16288 11933 16292
rect 11949 16348 12013 16352
rect 11949 16292 11953 16348
rect 11953 16292 12009 16348
rect 12009 16292 12013 16348
rect 11949 16288 12013 16292
rect 12029 16348 12093 16352
rect 12029 16292 12033 16348
rect 12033 16292 12089 16348
rect 12089 16292 12093 16348
rect 12029 16288 12093 16292
rect 12109 16348 12173 16352
rect 12109 16292 12113 16348
rect 12113 16292 12169 16348
rect 12169 16292 12173 16348
rect 12109 16288 12173 16292
rect 3681 15804 3745 15808
rect 3681 15748 3685 15804
rect 3685 15748 3741 15804
rect 3741 15748 3745 15804
rect 3681 15744 3745 15748
rect 3761 15804 3825 15808
rect 3761 15748 3765 15804
rect 3765 15748 3821 15804
rect 3821 15748 3825 15804
rect 3761 15744 3825 15748
rect 3841 15804 3905 15808
rect 3841 15748 3845 15804
rect 3845 15748 3901 15804
rect 3901 15748 3905 15804
rect 3841 15744 3905 15748
rect 3921 15804 3985 15808
rect 3921 15748 3925 15804
rect 3925 15748 3981 15804
rect 3981 15748 3985 15804
rect 3921 15744 3985 15748
rect 9140 15804 9204 15808
rect 9140 15748 9144 15804
rect 9144 15748 9200 15804
rect 9200 15748 9204 15804
rect 9140 15744 9204 15748
rect 9220 15804 9284 15808
rect 9220 15748 9224 15804
rect 9224 15748 9280 15804
rect 9280 15748 9284 15804
rect 9220 15744 9284 15748
rect 9300 15804 9364 15808
rect 9300 15748 9304 15804
rect 9304 15748 9360 15804
rect 9360 15748 9364 15804
rect 9300 15744 9364 15748
rect 9380 15804 9444 15808
rect 9380 15748 9384 15804
rect 9384 15748 9440 15804
rect 9440 15748 9444 15804
rect 9380 15744 9444 15748
rect 14598 15804 14662 15808
rect 14598 15748 14602 15804
rect 14602 15748 14658 15804
rect 14658 15748 14662 15804
rect 14598 15744 14662 15748
rect 14678 15804 14742 15808
rect 14678 15748 14682 15804
rect 14682 15748 14738 15804
rect 14738 15748 14742 15804
rect 14678 15744 14742 15748
rect 14758 15804 14822 15808
rect 14758 15748 14762 15804
rect 14762 15748 14818 15804
rect 14818 15748 14822 15804
rect 14758 15744 14822 15748
rect 14838 15804 14902 15808
rect 14838 15748 14842 15804
rect 14842 15748 14898 15804
rect 14898 15748 14902 15804
rect 14838 15744 14902 15748
rect 6410 15260 6474 15264
rect 6410 15204 6414 15260
rect 6414 15204 6470 15260
rect 6470 15204 6474 15260
rect 6410 15200 6474 15204
rect 6490 15260 6554 15264
rect 6490 15204 6494 15260
rect 6494 15204 6550 15260
rect 6550 15204 6554 15260
rect 6490 15200 6554 15204
rect 6570 15260 6634 15264
rect 6570 15204 6574 15260
rect 6574 15204 6630 15260
rect 6630 15204 6634 15260
rect 6570 15200 6634 15204
rect 6650 15260 6714 15264
rect 6650 15204 6654 15260
rect 6654 15204 6710 15260
rect 6710 15204 6714 15260
rect 6650 15200 6714 15204
rect 11869 15260 11933 15264
rect 11869 15204 11873 15260
rect 11873 15204 11929 15260
rect 11929 15204 11933 15260
rect 11869 15200 11933 15204
rect 11949 15260 12013 15264
rect 11949 15204 11953 15260
rect 11953 15204 12009 15260
rect 12009 15204 12013 15260
rect 11949 15200 12013 15204
rect 12029 15260 12093 15264
rect 12029 15204 12033 15260
rect 12033 15204 12089 15260
rect 12089 15204 12093 15260
rect 12029 15200 12093 15204
rect 12109 15260 12173 15264
rect 12109 15204 12113 15260
rect 12113 15204 12169 15260
rect 12169 15204 12173 15260
rect 12109 15200 12173 15204
rect 3681 14716 3745 14720
rect 3681 14660 3685 14716
rect 3685 14660 3741 14716
rect 3741 14660 3745 14716
rect 3681 14656 3745 14660
rect 3761 14716 3825 14720
rect 3761 14660 3765 14716
rect 3765 14660 3821 14716
rect 3821 14660 3825 14716
rect 3761 14656 3825 14660
rect 3841 14716 3905 14720
rect 3841 14660 3845 14716
rect 3845 14660 3901 14716
rect 3901 14660 3905 14716
rect 3841 14656 3905 14660
rect 3921 14716 3985 14720
rect 3921 14660 3925 14716
rect 3925 14660 3981 14716
rect 3981 14660 3985 14716
rect 3921 14656 3985 14660
rect 9140 14716 9204 14720
rect 9140 14660 9144 14716
rect 9144 14660 9200 14716
rect 9200 14660 9204 14716
rect 9140 14656 9204 14660
rect 9220 14716 9284 14720
rect 9220 14660 9224 14716
rect 9224 14660 9280 14716
rect 9280 14660 9284 14716
rect 9220 14656 9284 14660
rect 9300 14716 9364 14720
rect 9300 14660 9304 14716
rect 9304 14660 9360 14716
rect 9360 14660 9364 14716
rect 9300 14656 9364 14660
rect 9380 14716 9444 14720
rect 9380 14660 9384 14716
rect 9384 14660 9440 14716
rect 9440 14660 9444 14716
rect 9380 14656 9444 14660
rect 14598 14716 14662 14720
rect 14598 14660 14602 14716
rect 14602 14660 14658 14716
rect 14658 14660 14662 14716
rect 14598 14656 14662 14660
rect 14678 14716 14742 14720
rect 14678 14660 14682 14716
rect 14682 14660 14738 14716
rect 14738 14660 14742 14716
rect 14678 14656 14742 14660
rect 14758 14716 14822 14720
rect 14758 14660 14762 14716
rect 14762 14660 14818 14716
rect 14818 14660 14822 14716
rect 14758 14656 14822 14660
rect 14838 14716 14902 14720
rect 14838 14660 14842 14716
rect 14842 14660 14898 14716
rect 14898 14660 14902 14716
rect 14838 14656 14902 14660
rect 6410 14172 6474 14176
rect 6410 14116 6414 14172
rect 6414 14116 6470 14172
rect 6470 14116 6474 14172
rect 6410 14112 6474 14116
rect 6490 14172 6554 14176
rect 6490 14116 6494 14172
rect 6494 14116 6550 14172
rect 6550 14116 6554 14172
rect 6490 14112 6554 14116
rect 6570 14172 6634 14176
rect 6570 14116 6574 14172
rect 6574 14116 6630 14172
rect 6630 14116 6634 14172
rect 6570 14112 6634 14116
rect 6650 14172 6714 14176
rect 6650 14116 6654 14172
rect 6654 14116 6710 14172
rect 6710 14116 6714 14172
rect 6650 14112 6714 14116
rect 11869 14172 11933 14176
rect 11869 14116 11873 14172
rect 11873 14116 11929 14172
rect 11929 14116 11933 14172
rect 11869 14112 11933 14116
rect 11949 14172 12013 14176
rect 11949 14116 11953 14172
rect 11953 14116 12009 14172
rect 12009 14116 12013 14172
rect 11949 14112 12013 14116
rect 12029 14172 12093 14176
rect 12029 14116 12033 14172
rect 12033 14116 12089 14172
rect 12089 14116 12093 14172
rect 12029 14112 12093 14116
rect 12109 14172 12173 14176
rect 12109 14116 12113 14172
rect 12113 14116 12169 14172
rect 12169 14116 12173 14172
rect 12109 14112 12173 14116
rect 3681 13628 3745 13632
rect 3681 13572 3685 13628
rect 3685 13572 3741 13628
rect 3741 13572 3745 13628
rect 3681 13568 3745 13572
rect 3761 13628 3825 13632
rect 3761 13572 3765 13628
rect 3765 13572 3821 13628
rect 3821 13572 3825 13628
rect 3761 13568 3825 13572
rect 3841 13628 3905 13632
rect 3841 13572 3845 13628
rect 3845 13572 3901 13628
rect 3901 13572 3905 13628
rect 3841 13568 3905 13572
rect 3921 13628 3985 13632
rect 3921 13572 3925 13628
rect 3925 13572 3981 13628
rect 3981 13572 3985 13628
rect 3921 13568 3985 13572
rect 9140 13628 9204 13632
rect 9140 13572 9144 13628
rect 9144 13572 9200 13628
rect 9200 13572 9204 13628
rect 9140 13568 9204 13572
rect 9220 13628 9284 13632
rect 9220 13572 9224 13628
rect 9224 13572 9280 13628
rect 9280 13572 9284 13628
rect 9220 13568 9284 13572
rect 9300 13628 9364 13632
rect 9300 13572 9304 13628
rect 9304 13572 9360 13628
rect 9360 13572 9364 13628
rect 9300 13568 9364 13572
rect 9380 13628 9444 13632
rect 9380 13572 9384 13628
rect 9384 13572 9440 13628
rect 9440 13572 9444 13628
rect 9380 13568 9444 13572
rect 14598 13628 14662 13632
rect 14598 13572 14602 13628
rect 14602 13572 14658 13628
rect 14658 13572 14662 13628
rect 14598 13568 14662 13572
rect 14678 13628 14742 13632
rect 14678 13572 14682 13628
rect 14682 13572 14738 13628
rect 14738 13572 14742 13628
rect 14678 13568 14742 13572
rect 14758 13628 14822 13632
rect 14758 13572 14762 13628
rect 14762 13572 14818 13628
rect 14818 13572 14822 13628
rect 14758 13568 14822 13572
rect 14838 13628 14902 13632
rect 14838 13572 14842 13628
rect 14842 13572 14898 13628
rect 14898 13572 14902 13628
rect 14838 13568 14902 13572
rect 6410 13084 6474 13088
rect 6410 13028 6414 13084
rect 6414 13028 6470 13084
rect 6470 13028 6474 13084
rect 6410 13024 6474 13028
rect 6490 13084 6554 13088
rect 6490 13028 6494 13084
rect 6494 13028 6550 13084
rect 6550 13028 6554 13084
rect 6490 13024 6554 13028
rect 6570 13084 6634 13088
rect 6570 13028 6574 13084
rect 6574 13028 6630 13084
rect 6630 13028 6634 13084
rect 6570 13024 6634 13028
rect 6650 13084 6714 13088
rect 6650 13028 6654 13084
rect 6654 13028 6710 13084
rect 6710 13028 6714 13084
rect 6650 13024 6714 13028
rect 11869 13084 11933 13088
rect 11869 13028 11873 13084
rect 11873 13028 11929 13084
rect 11929 13028 11933 13084
rect 11869 13024 11933 13028
rect 11949 13084 12013 13088
rect 11949 13028 11953 13084
rect 11953 13028 12009 13084
rect 12009 13028 12013 13084
rect 11949 13024 12013 13028
rect 12029 13084 12093 13088
rect 12029 13028 12033 13084
rect 12033 13028 12089 13084
rect 12089 13028 12093 13084
rect 12029 13024 12093 13028
rect 12109 13084 12173 13088
rect 12109 13028 12113 13084
rect 12113 13028 12169 13084
rect 12169 13028 12173 13084
rect 12109 13024 12173 13028
rect 3681 12540 3745 12544
rect 3681 12484 3685 12540
rect 3685 12484 3741 12540
rect 3741 12484 3745 12540
rect 3681 12480 3745 12484
rect 3761 12540 3825 12544
rect 3761 12484 3765 12540
rect 3765 12484 3821 12540
rect 3821 12484 3825 12540
rect 3761 12480 3825 12484
rect 3841 12540 3905 12544
rect 3841 12484 3845 12540
rect 3845 12484 3901 12540
rect 3901 12484 3905 12540
rect 3841 12480 3905 12484
rect 3921 12540 3985 12544
rect 3921 12484 3925 12540
rect 3925 12484 3981 12540
rect 3981 12484 3985 12540
rect 3921 12480 3985 12484
rect 9140 12540 9204 12544
rect 9140 12484 9144 12540
rect 9144 12484 9200 12540
rect 9200 12484 9204 12540
rect 9140 12480 9204 12484
rect 9220 12540 9284 12544
rect 9220 12484 9224 12540
rect 9224 12484 9280 12540
rect 9280 12484 9284 12540
rect 9220 12480 9284 12484
rect 9300 12540 9364 12544
rect 9300 12484 9304 12540
rect 9304 12484 9360 12540
rect 9360 12484 9364 12540
rect 9300 12480 9364 12484
rect 9380 12540 9444 12544
rect 9380 12484 9384 12540
rect 9384 12484 9440 12540
rect 9440 12484 9444 12540
rect 9380 12480 9444 12484
rect 14598 12540 14662 12544
rect 14598 12484 14602 12540
rect 14602 12484 14658 12540
rect 14658 12484 14662 12540
rect 14598 12480 14662 12484
rect 14678 12540 14742 12544
rect 14678 12484 14682 12540
rect 14682 12484 14738 12540
rect 14738 12484 14742 12540
rect 14678 12480 14742 12484
rect 14758 12540 14822 12544
rect 14758 12484 14762 12540
rect 14762 12484 14818 12540
rect 14818 12484 14822 12540
rect 14758 12480 14822 12484
rect 14838 12540 14902 12544
rect 14838 12484 14842 12540
rect 14842 12484 14898 12540
rect 14898 12484 14902 12540
rect 14838 12480 14902 12484
rect 6410 11996 6474 12000
rect 6410 11940 6414 11996
rect 6414 11940 6470 11996
rect 6470 11940 6474 11996
rect 6410 11936 6474 11940
rect 6490 11996 6554 12000
rect 6490 11940 6494 11996
rect 6494 11940 6550 11996
rect 6550 11940 6554 11996
rect 6490 11936 6554 11940
rect 6570 11996 6634 12000
rect 6570 11940 6574 11996
rect 6574 11940 6630 11996
rect 6630 11940 6634 11996
rect 6570 11936 6634 11940
rect 6650 11996 6714 12000
rect 6650 11940 6654 11996
rect 6654 11940 6710 11996
rect 6710 11940 6714 11996
rect 6650 11936 6714 11940
rect 11869 11996 11933 12000
rect 11869 11940 11873 11996
rect 11873 11940 11929 11996
rect 11929 11940 11933 11996
rect 11869 11936 11933 11940
rect 11949 11996 12013 12000
rect 11949 11940 11953 11996
rect 11953 11940 12009 11996
rect 12009 11940 12013 11996
rect 11949 11936 12013 11940
rect 12029 11996 12093 12000
rect 12029 11940 12033 11996
rect 12033 11940 12089 11996
rect 12089 11940 12093 11996
rect 12029 11936 12093 11940
rect 12109 11996 12173 12000
rect 12109 11940 12113 11996
rect 12113 11940 12169 11996
rect 12169 11940 12173 11996
rect 12109 11936 12173 11940
rect 3681 11452 3745 11456
rect 3681 11396 3685 11452
rect 3685 11396 3741 11452
rect 3741 11396 3745 11452
rect 3681 11392 3745 11396
rect 3761 11452 3825 11456
rect 3761 11396 3765 11452
rect 3765 11396 3821 11452
rect 3821 11396 3825 11452
rect 3761 11392 3825 11396
rect 3841 11452 3905 11456
rect 3841 11396 3845 11452
rect 3845 11396 3901 11452
rect 3901 11396 3905 11452
rect 3841 11392 3905 11396
rect 3921 11452 3985 11456
rect 3921 11396 3925 11452
rect 3925 11396 3981 11452
rect 3981 11396 3985 11452
rect 3921 11392 3985 11396
rect 9140 11452 9204 11456
rect 9140 11396 9144 11452
rect 9144 11396 9200 11452
rect 9200 11396 9204 11452
rect 9140 11392 9204 11396
rect 9220 11452 9284 11456
rect 9220 11396 9224 11452
rect 9224 11396 9280 11452
rect 9280 11396 9284 11452
rect 9220 11392 9284 11396
rect 9300 11452 9364 11456
rect 9300 11396 9304 11452
rect 9304 11396 9360 11452
rect 9360 11396 9364 11452
rect 9300 11392 9364 11396
rect 9380 11452 9444 11456
rect 9380 11396 9384 11452
rect 9384 11396 9440 11452
rect 9440 11396 9444 11452
rect 9380 11392 9444 11396
rect 14598 11452 14662 11456
rect 14598 11396 14602 11452
rect 14602 11396 14658 11452
rect 14658 11396 14662 11452
rect 14598 11392 14662 11396
rect 14678 11452 14742 11456
rect 14678 11396 14682 11452
rect 14682 11396 14738 11452
rect 14738 11396 14742 11452
rect 14678 11392 14742 11396
rect 14758 11452 14822 11456
rect 14758 11396 14762 11452
rect 14762 11396 14818 11452
rect 14818 11396 14822 11452
rect 14758 11392 14822 11396
rect 14838 11452 14902 11456
rect 14838 11396 14842 11452
rect 14842 11396 14898 11452
rect 14898 11396 14902 11452
rect 14838 11392 14902 11396
rect 6410 10908 6474 10912
rect 6410 10852 6414 10908
rect 6414 10852 6470 10908
rect 6470 10852 6474 10908
rect 6410 10848 6474 10852
rect 6490 10908 6554 10912
rect 6490 10852 6494 10908
rect 6494 10852 6550 10908
rect 6550 10852 6554 10908
rect 6490 10848 6554 10852
rect 6570 10908 6634 10912
rect 6570 10852 6574 10908
rect 6574 10852 6630 10908
rect 6630 10852 6634 10908
rect 6570 10848 6634 10852
rect 6650 10908 6714 10912
rect 6650 10852 6654 10908
rect 6654 10852 6710 10908
rect 6710 10852 6714 10908
rect 6650 10848 6714 10852
rect 11869 10908 11933 10912
rect 11869 10852 11873 10908
rect 11873 10852 11929 10908
rect 11929 10852 11933 10908
rect 11869 10848 11933 10852
rect 11949 10908 12013 10912
rect 11949 10852 11953 10908
rect 11953 10852 12009 10908
rect 12009 10852 12013 10908
rect 11949 10848 12013 10852
rect 12029 10908 12093 10912
rect 12029 10852 12033 10908
rect 12033 10852 12089 10908
rect 12089 10852 12093 10908
rect 12029 10848 12093 10852
rect 12109 10908 12173 10912
rect 12109 10852 12113 10908
rect 12113 10852 12169 10908
rect 12169 10852 12173 10908
rect 12109 10848 12173 10852
rect 3681 10364 3745 10368
rect 3681 10308 3685 10364
rect 3685 10308 3741 10364
rect 3741 10308 3745 10364
rect 3681 10304 3745 10308
rect 3761 10364 3825 10368
rect 3761 10308 3765 10364
rect 3765 10308 3821 10364
rect 3821 10308 3825 10364
rect 3761 10304 3825 10308
rect 3841 10364 3905 10368
rect 3841 10308 3845 10364
rect 3845 10308 3901 10364
rect 3901 10308 3905 10364
rect 3841 10304 3905 10308
rect 3921 10364 3985 10368
rect 3921 10308 3925 10364
rect 3925 10308 3981 10364
rect 3981 10308 3985 10364
rect 3921 10304 3985 10308
rect 9140 10364 9204 10368
rect 9140 10308 9144 10364
rect 9144 10308 9200 10364
rect 9200 10308 9204 10364
rect 9140 10304 9204 10308
rect 9220 10364 9284 10368
rect 9220 10308 9224 10364
rect 9224 10308 9280 10364
rect 9280 10308 9284 10364
rect 9220 10304 9284 10308
rect 9300 10364 9364 10368
rect 9300 10308 9304 10364
rect 9304 10308 9360 10364
rect 9360 10308 9364 10364
rect 9300 10304 9364 10308
rect 9380 10364 9444 10368
rect 9380 10308 9384 10364
rect 9384 10308 9440 10364
rect 9440 10308 9444 10364
rect 9380 10304 9444 10308
rect 14598 10364 14662 10368
rect 14598 10308 14602 10364
rect 14602 10308 14658 10364
rect 14658 10308 14662 10364
rect 14598 10304 14662 10308
rect 14678 10364 14742 10368
rect 14678 10308 14682 10364
rect 14682 10308 14738 10364
rect 14738 10308 14742 10364
rect 14678 10304 14742 10308
rect 14758 10364 14822 10368
rect 14758 10308 14762 10364
rect 14762 10308 14818 10364
rect 14818 10308 14822 10364
rect 14758 10304 14822 10308
rect 14838 10364 14902 10368
rect 14838 10308 14842 10364
rect 14842 10308 14898 10364
rect 14898 10308 14902 10364
rect 14838 10304 14902 10308
rect 6410 9820 6474 9824
rect 6410 9764 6414 9820
rect 6414 9764 6470 9820
rect 6470 9764 6474 9820
rect 6410 9760 6474 9764
rect 6490 9820 6554 9824
rect 6490 9764 6494 9820
rect 6494 9764 6550 9820
rect 6550 9764 6554 9820
rect 6490 9760 6554 9764
rect 6570 9820 6634 9824
rect 6570 9764 6574 9820
rect 6574 9764 6630 9820
rect 6630 9764 6634 9820
rect 6570 9760 6634 9764
rect 6650 9820 6714 9824
rect 6650 9764 6654 9820
rect 6654 9764 6710 9820
rect 6710 9764 6714 9820
rect 6650 9760 6714 9764
rect 11869 9820 11933 9824
rect 11869 9764 11873 9820
rect 11873 9764 11929 9820
rect 11929 9764 11933 9820
rect 11869 9760 11933 9764
rect 11949 9820 12013 9824
rect 11949 9764 11953 9820
rect 11953 9764 12009 9820
rect 12009 9764 12013 9820
rect 11949 9760 12013 9764
rect 12029 9820 12093 9824
rect 12029 9764 12033 9820
rect 12033 9764 12089 9820
rect 12089 9764 12093 9820
rect 12029 9760 12093 9764
rect 12109 9820 12173 9824
rect 12109 9764 12113 9820
rect 12113 9764 12169 9820
rect 12169 9764 12173 9820
rect 12109 9760 12173 9764
rect 3681 9276 3745 9280
rect 3681 9220 3685 9276
rect 3685 9220 3741 9276
rect 3741 9220 3745 9276
rect 3681 9216 3745 9220
rect 3761 9276 3825 9280
rect 3761 9220 3765 9276
rect 3765 9220 3821 9276
rect 3821 9220 3825 9276
rect 3761 9216 3825 9220
rect 3841 9276 3905 9280
rect 3841 9220 3845 9276
rect 3845 9220 3901 9276
rect 3901 9220 3905 9276
rect 3841 9216 3905 9220
rect 3921 9276 3985 9280
rect 3921 9220 3925 9276
rect 3925 9220 3981 9276
rect 3981 9220 3985 9276
rect 3921 9216 3985 9220
rect 9140 9276 9204 9280
rect 9140 9220 9144 9276
rect 9144 9220 9200 9276
rect 9200 9220 9204 9276
rect 9140 9216 9204 9220
rect 9220 9276 9284 9280
rect 9220 9220 9224 9276
rect 9224 9220 9280 9276
rect 9280 9220 9284 9276
rect 9220 9216 9284 9220
rect 9300 9276 9364 9280
rect 9300 9220 9304 9276
rect 9304 9220 9360 9276
rect 9360 9220 9364 9276
rect 9300 9216 9364 9220
rect 9380 9276 9444 9280
rect 9380 9220 9384 9276
rect 9384 9220 9440 9276
rect 9440 9220 9444 9276
rect 9380 9216 9444 9220
rect 14598 9276 14662 9280
rect 14598 9220 14602 9276
rect 14602 9220 14658 9276
rect 14658 9220 14662 9276
rect 14598 9216 14662 9220
rect 14678 9276 14742 9280
rect 14678 9220 14682 9276
rect 14682 9220 14738 9276
rect 14738 9220 14742 9276
rect 14678 9216 14742 9220
rect 14758 9276 14822 9280
rect 14758 9220 14762 9276
rect 14762 9220 14818 9276
rect 14818 9220 14822 9276
rect 14758 9216 14822 9220
rect 14838 9276 14902 9280
rect 14838 9220 14842 9276
rect 14842 9220 14898 9276
rect 14898 9220 14902 9276
rect 14838 9216 14902 9220
rect 6410 8732 6474 8736
rect 6410 8676 6414 8732
rect 6414 8676 6470 8732
rect 6470 8676 6474 8732
rect 6410 8672 6474 8676
rect 6490 8732 6554 8736
rect 6490 8676 6494 8732
rect 6494 8676 6550 8732
rect 6550 8676 6554 8732
rect 6490 8672 6554 8676
rect 6570 8732 6634 8736
rect 6570 8676 6574 8732
rect 6574 8676 6630 8732
rect 6630 8676 6634 8732
rect 6570 8672 6634 8676
rect 6650 8732 6714 8736
rect 6650 8676 6654 8732
rect 6654 8676 6710 8732
rect 6710 8676 6714 8732
rect 6650 8672 6714 8676
rect 11869 8732 11933 8736
rect 11869 8676 11873 8732
rect 11873 8676 11929 8732
rect 11929 8676 11933 8732
rect 11869 8672 11933 8676
rect 11949 8732 12013 8736
rect 11949 8676 11953 8732
rect 11953 8676 12009 8732
rect 12009 8676 12013 8732
rect 11949 8672 12013 8676
rect 12029 8732 12093 8736
rect 12029 8676 12033 8732
rect 12033 8676 12089 8732
rect 12089 8676 12093 8732
rect 12029 8672 12093 8676
rect 12109 8732 12173 8736
rect 12109 8676 12113 8732
rect 12113 8676 12169 8732
rect 12169 8676 12173 8732
rect 12109 8672 12173 8676
rect 3681 8188 3745 8192
rect 3681 8132 3685 8188
rect 3685 8132 3741 8188
rect 3741 8132 3745 8188
rect 3681 8128 3745 8132
rect 3761 8188 3825 8192
rect 3761 8132 3765 8188
rect 3765 8132 3821 8188
rect 3821 8132 3825 8188
rect 3761 8128 3825 8132
rect 3841 8188 3905 8192
rect 3841 8132 3845 8188
rect 3845 8132 3901 8188
rect 3901 8132 3905 8188
rect 3841 8128 3905 8132
rect 3921 8188 3985 8192
rect 3921 8132 3925 8188
rect 3925 8132 3981 8188
rect 3981 8132 3985 8188
rect 3921 8128 3985 8132
rect 9140 8188 9204 8192
rect 9140 8132 9144 8188
rect 9144 8132 9200 8188
rect 9200 8132 9204 8188
rect 9140 8128 9204 8132
rect 9220 8188 9284 8192
rect 9220 8132 9224 8188
rect 9224 8132 9280 8188
rect 9280 8132 9284 8188
rect 9220 8128 9284 8132
rect 9300 8188 9364 8192
rect 9300 8132 9304 8188
rect 9304 8132 9360 8188
rect 9360 8132 9364 8188
rect 9300 8128 9364 8132
rect 9380 8188 9444 8192
rect 9380 8132 9384 8188
rect 9384 8132 9440 8188
rect 9440 8132 9444 8188
rect 9380 8128 9444 8132
rect 14598 8188 14662 8192
rect 14598 8132 14602 8188
rect 14602 8132 14658 8188
rect 14658 8132 14662 8188
rect 14598 8128 14662 8132
rect 14678 8188 14742 8192
rect 14678 8132 14682 8188
rect 14682 8132 14738 8188
rect 14738 8132 14742 8188
rect 14678 8128 14742 8132
rect 14758 8188 14822 8192
rect 14758 8132 14762 8188
rect 14762 8132 14818 8188
rect 14818 8132 14822 8188
rect 14758 8128 14822 8132
rect 14838 8188 14902 8192
rect 14838 8132 14842 8188
rect 14842 8132 14898 8188
rect 14898 8132 14902 8188
rect 14838 8128 14902 8132
rect 6410 7644 6474 7648
rect 6410 7588 6414 7644
rect 6414 7588 6470 7644
rect 6470 7588 6474 7644
rect 6410 7584 6474 7588
rect 6490 7644 6554 7648
rect 6490 7588 6494 7644
rect 6494 7588 6550 7644
rect 6550 7588 6554 7644
rect 6490 7584 6554 7588
rect 6570 7644 6634 7648
rect 6570 7588 6574 7644
rect 6574 7588 6630 7644
rect 6630 7588 6634 7644
rect 6570 7584 6634 7588
rect 6650 7644 6714 7648
rect 6650 7588 6654 7644
rect 6654 7588 6710 7644
rect 6710 7588 6714 7644
rect 6650 7584 6714 7588
rect 11869 7644 11933 7648
rect 11869 7588 11873 7644
rect 11873 7588 11929 7644
rect 11929 7588 11933 7644
rect 11869 7584 11933 7588
rect 11949 7644 12013 7648
rect 11949 7588 11953 7644
rect 11953 7588 12009 7644
rect 12009 7588 12013 7644
rect 11949 7584 12013 7588
rect 12029 7644 12093 7648
rect 12029 7588 12033 7644
rect 12033 7588 12089 7644
rect 12089 7588 12093 7644
rect 12029 7584 12093 7588
rect 12109 7644 12173 7648
rect 12109 7588 12113 7644
rect 12113 7588 12169 7644
rect 12169 7588 12173 7644
rect 12109 7584 12173 7588
rect 3681 7100 3745 7104
rect 3681 7044 3685 7100
rect 3685 7044 3741 7100
rect 3741 7044 3745 7100
rect 3681 7040 3745 7044
rect 3761 7100 3825 7104
rect 3761 7044 3765 7100
rect 3765 7044 3821 7100
rect 3821 7044 3825 7100
rect 3761 7040 3825 7044
rect 3841 7100 3905 7104
rect 3841 7044 3845 7100
rect 3845 7044 3901 7100
rect 3901 7044 3905 7100
rect 3841 7040 3905 7044
rect 3921 7100 3985 7104
rect 3921 7044 3925 7100
rect 3925 7044 3981 7100
rect 3981 7044 3985 7100
rect 3921 7040 3985 7044
rect 9140 7100 9204 7104
rect 9140 7044 9144 7100
rect 9144 7044 9200 7100
rect 9200 7044 9204 7100
rect 9140 7040 9204 7044
rect 9220 7100 9284 7104
rect 9220 7044 9224 7100
rect 9224 7044 9280 7100
rect 9280 7044 9284 7100
rect 9220 7040 9284 7044
rect 9300 7100 9364 7104
rect 9300 7044 9304 7100
rect 9304 7044 9360 7100
rect 9360 7044 9364 7100
rect 9300 7040 9364 7044
rect 9380 7100 9444 7104
rect 9380 7044 9384 7100
rect 9384 7044 9440 7100
rect 9440 7044 9444 7100
rect 9380 7040 9444 7044
rect 14598 7100 14662 7104
rect 14598 7044 14602 7100
rect 14602 7044 14658 7100
rect 14658 7044 14662 7100
rect 14598 7040 14662 7044
rect 14678 7100 14742 7104
rect 14678 7044 14682 7100
rect 14682 7044 14738 7100
rect 14738 7044 14742 7100
rect 14678 7040 14742 7044
rect 14758 7100 14822 7104
rect 14758 7044 14762 7100
rect 14762 7044 14818 7100
rect 14818 7044 14822 7100
rect 14758 7040 14822 7044
rect 14838 7100 14902 7104
rect 14838 7044 14842 7100
rect 14842 7044 14898 7100
rect 14898 7044 14902 7100
rect 14838 7040 14902 7044
rect 6410 6556 6474 6560
rect 6410 6500 6414 6556
rect 6414 6500 6470 6556
rect 6470 6500 6474 6556
rect 6410 6496 6474 6500
rect 6490 6556 6554 6560
rect 6490 6500 6494 6556
rect 6494 6500 6550 6556
rect 6550 6500 6554 6556
rect 6490 6496 6554 6500
rect 6570 6556 6634 6560
rect 6570 6500 6574 6556
rect 6574 6500 6630 6556
rect 6630 6500 6634 6556
rect 6570 6496 6634 6500
rect 6650 6556 6714 6560
rect 6650 6500 6654 6556
rect 6654 6500 6710 6556
rect 6710 6500 6714 6556
rect 6650 6496 6714 6500
rect 11869 6556 11933 6560
rect 11869 6500 11873 6556
rect 11873 6500 11929 6556
rect 11929 6500 11933 6556
rect 11869 6496 11933 6500
rect 11949 6556 12013 6560
rect 11949 6500 11953 6556
rect 11953 6500 12009 6556
rect 12009 6500 12013 6556
rect 11949 6496 12013 6500
rect 12029 6556 12093 6560
rect 12029 6500 12033 6556
rect 12033 6500 12089 6556
rect 12089 6500 12093 6556
rect 12029 6496 12093 6500
rect 12109 6556 12173 6560
rect 12109 6500 12113 6556
rect 12113 6500 12169 6556
rect 12169 6500 12173 6556
rect 12109 6496 12173 6500
rect 3681 6012 3745 6016
rect 3681 5956 3685 6012
rect 3685 5956 3741 6012
rect 3741 5956 3745 6012
rect 3681 5952 3745 5956
rect 3761 6012 3825 6016
rect 3761 5956 3765 6012
rect 3765 5956 3821 6012
rect 3821 5956 3825 6012
rect 3761 5952 3825 5956
rect 3841 6012 3905 6016
rect 3841 5956 3845 6012
rect 3845 5956 3901 6012
rect 3901 5956 3905 6012
rect 3841 5952 3905 5956
rect 3921 6012 3985 6016
rect 3921 5956 3925 6012
rect 3925 5956 3981 6012
rect 3981 5956 3985 6012
rect 3921 5952 3985 5956
rect 9140 6012 9204 6016
rect 9140 5956 9144 6012
rect 9144 5956 9200 6012
rect 9200 5956 9204 6012
rect 9140 5952 9204 5956
rect 9220 6012 9284 6016
rect 9220 5956 9224 6012
rect 9224 5956 9280 6012
rect 9280 5956 9284 6012
rect 9220 5952 9284 5956
rect 9300 6012 9364 6016
rect 9300 5956 9304 6012
rect 9304 5956 9360 6012
rect 9360 5956 9364 6012
rect 9300 5952 9364 5956
rect 9380 6012 9444 6016
rect 9380 5956 9384 6012
rect 9384 5956 9440 6012
rect 9440 5956 9444 6012
rect 9380 5952 9444 5956
rect 14598 6012 14662 6016
rect 14598 5956 14602 6012
rect 14602 5956 14658 6012
rect 14658 5956 14662 6012
rect 14598 5952 14662 5956
rect 14678 6012 14742 6016
rect 14678 5956 14682 6012
rect 14682 5956 14738 6012
rect 14738 5956 14742 6012
rect 14678 5952 14742 5956
rect 14758 6012 14822 6016
rect 14758 5956 14762 6012
rect 14762 5956 14818 6012
rect 14818 5956 14822 6012
rect 14758 5952 14822 5956
rect 14838 6012 14902 6016
rect 14838 5956 14842 6012
rect 14842 5956 14898 6012
rect 14898 5956 14902 6012
rect 14838 5952 14902 5956
rect 6410 5468 6474 5472
rect 6410 5412 6414 5468
rect 6414 5412 6470 5468
rect 6470 5412 6474 5468
rect 6410 5408 6474 5412
rect 6490 5468 6554 5472
rect 6490 5412 6494 5468
rect 6494 5412 6550 5468
rect 6550 5412 6554 5468
rect 6490 5408 6554 5412
rect 6570 5468 6634 5472
rect 6570 5412 6574 5468
rect 6574 5412 6630 5468
rect 6630 5412 6634 5468
rect 6570 5408 6634 5412
rect 6650 5468 6714 5472
rect 6650 5412 6654 5468
rect 6654 5412 6710 5468
rect 6710 5412 6714 5468
rect 6650 5408 6714 5412
rect 11869 5468 11933 5472
rect 11869 5412 11873 5468
rect 11873 5412 11929 5468
rect 11929 5412 11933 5468
rect 11869 5408 11933 5412
rect 11949 5468 12013 5472
rect 11949 5412 11953 5468
rect 11953 5412 12009 5468
rect 12009 5412 12013 5468
rect 11949 5408 12013 5412
rect 12029 5468 12093 5472
rect 12029 5412 12033 5468
rect 12033 5412 12089 5468
rect 12089 5412 12093 5468
rect 12029 5408 12093 5412
rect 12109 5468 12173 5472
rect 12109 5412 12113 5468
rect 12113 5412 12169 5468
rect 12169 5412 12173 5468
rect 12109 5408 12173 5412
rect 3681 4924 3745 4928
rect 3681 4868 3685 4924
rect 3685 4868 3741 4924
rect 3741 4868 3745 4924
rect 3681 4864 3745 4868
rect 3761 4924 3825 4928
rect 3761 4868 3765 4924
rect 3765 4868 3821 4924
rect 3821 4868 3825 4924
rect 3761 4864 3825 4868
rect 3841 4924 3905 4928
rect 3841 4868 3845 4924
rect 3845 4868 3901 4924
rect 3901 4868 3905 4924
rect 3841 4864 3905 4868
rect 3921 4924 3985 4928
rect 3921 4868 3925 4924
rect 3925 4868 3981 4924
rect 3981 4868 3985 4924
rect 3921 4864 3985 4868
rect 9140 4924 9204 4928
rect 9140 4868 9144 4924
rect 9144 4868 9200 4924
rect 9200 4868 9204 4924
rect 9140 4864 9204 4868
rect 9220 4924 9284 4928
rect 9220 4868 9224 4924
rect 9224 4868 9280 4924
rect 9280 4868 9284 4924
rect 9220 4864 9284 4868
rect 9300 4924 9364 4928
rect 9300 4868 9304 4924
rect 9304 4868 9360 4924
rect 9360 4868 9364 4924
rect 9300 4864 9364 4868
rect 9380 4924 9444 4928
rect 9380 4868 9384 4924
rect 9384 4868 9440 4924
rect 9440 4868 9444 4924
rect 9380 4864 9444 4868
rect 14598 4924 14662 4928
rect 14598 4868 14602 4924
rect 14602 4868 14658 4924
rect 14658 4868 14662 4924
rect 14598 4864 14662 4868
rect 14678 4924 14742 4928
rect 14678 4868 14682 4924
rect 14682 4868 14738 4924
rect 14738 4868 14742 4924
rect 14678 4864 14742 4868
rect 14758 4924 14822 4928
rect 14758 4868 14762 4924
rect 14762 4868 14818 4924
rect 14818 4868 14822 4924
rect 14758 4864 14822 4868
rect 14838 4924 14902 4928
rect 14838 4868 14842 4924
rect 14842 4868 14898 4924
rect 14898 4868 14902 4924
rect 14838 4864 14902 4868
rect 6410 4380 6474 4384
rect 6410 4324 6414 4380
rect 6414 4324 6470 4380
rect 6470 4324 6474 4380
rect 6410 4320 6474 4324
rect 6490 4380 6554 4384
rect 6490 4324 6494 4380
rect 6494 4324 6550 4380
rect 6550 4324 6554 4380
rect 6490 4320 6554 4324
rect 6570 4380 6634 4384
rect 6570 4324 6574 4380
rect 6574 4324 6630 4380
rect 6630 4324 6634 4380
rect 6570 4320 6634 4324
rect 6650 4380 6714 4384
rect 6650 4324 6654 4380
rect 6654 4324 6710 4380
rect 6710 4324 6714 4380
rect 6650 4320 6714 4324
rect 11869 4380 11933 4384
rect 11869 4324 11873 4380
rect 11873 4324 11929 4380
rect 11929 4324 11933 4380
rect 11869 4320 11933 4324
rect 11949 4380 12013 4384
rect 11949 4324 11953 4380
rect 11953 4324 12009 4380
rect 12009 4324 12013 4380
rect 11949 4320 12013 4324
rect 12029 4380 12093 4384
rect 12029 4324 12033 4380
rect 12033 4324 12089 4380
rect 12089 4324 12093 4380
rect 12029 4320 12093 4324
rect 12109 4380 12173 4384
rect 12109 4324 12113 4380
rect 12113 4324 12169 4380
rect 12169 4324 12173 4380
rect 12109 4320 12173 4324
rect 3681 3836 3745 3840
rect 3681 3780 3685 3836
rect 3685 3780 3741 3836
rect 3741 3780 3745 3836
rect 3681 3776 3745 3780
rect 3761 3836 3825 3840
rect 3761 3780 3765 3836
rect 3765 3780 3821 3836
rect 3821 3780 3825 3836
rect 3761 3776 3825 3780
rect 3841 3836 3905 3840
rect 3841 3780 3845 3836
rect 3845 3780 3901 3836
rect 3901 3780 3905 3836
rect 3841 3776 3905 3780
rect 3921 3836 3985 3840
rect 3921 3780 3925 3836
rect 3925 3780 3981 3836
rect 3981 3780 3985 3836
rect 3921 3776 3985 3780
rect 9140 3836 9204 3840
rect 9140 3780 9144 3836
rect 9144 3780 9200 3836
rect 9200 3780 9204 3836
rect 9140 3776 9204 3780
rect 9220 3836 9284 3840
rect 9220 3780 9224 3836
rect 9224 3780 9280 3836
rect 9280 3780 9284 3836
rect 9220 3776 9284 3780
rect 9300 3836 9364 3840
rect 9300 3780 9304 3836
rect 9304 3780 9360 3836
rect 9360 3780 9364 3836
rect 9300 3776 9364 3780
rect 9380 3836 9444 3840
rect 9380 3780 9384 3836
rect 9384 3780 9440 3836
rect 9440 3780 9444 3836
rect 9380 3776 9444 3780
rect 14598 3836 14662 3840
rect 14598 3780 14602 3836
rect 14602 3780 14658 3836
rect 14658 3780 14662 3836
rect 14598 3776 14662 3780
rect 14678 3836 14742 3840
rect 14678 3780 14682 3836
rect 14682 3780 14738 3836
rect 14738 3780 14742 3836
rect 14678 3776 14742 3780
rect 14758 3836 14822 3840
rect 14758 3780 14762 3836
rect 14762 3780 14818 3836
rect 14818 3780 14822 3836
rect 14758 3776 14822 3780
rect 14838 3836 14902 3840
rect 14838 3780 14842 3836
rect 14842 3780 14898 3836
rect 14898 3780 14902 3836
rect 14838 3776 14902 3780
rect 6410 3292 6474 3296
rect 6410 3236 6414 3292
rect 6414 3236 6470 3292
rect 6470 3236 6474 3292
rect 6410 3232 6474 3236
rect 6490 3292 6554 3296
rect 6490 3236 6494 3292
rect 6494 3236 6550 3292
rect 6550 3236 6554 3292
rect 6490 3232 6554 3236
rect 6570 3292 6634 3296
rect 6570 3236 6574 3292
rect 6574 3236 6630 3292
rect 6630 3236 6634 3292
rect 6570 3232 6634 3236
rect 6650 3292 6714 3296
rect 6650 3236 6654 3292
rect 6654 3236 6710 3292
rect 6710 3236 6714 3292
rect 6650 3232 6714 3236
rect 11869 3292 11933 3296
rect 11869 3236 11873 3292
rect 11873 3236 11929 3292
rect 11929 3236 11933 3292
rect 11869 3232 11933 3236
rect 11949 3292 12013 3296
rect 11949 3236 11953 3292
rect 11953 3236 12009 3292
rect 12009 3236 12013 3292
rect 11949 3232 12013 3236
rect 12029 3292 12093 3296
rect 12029 3236 12033 3292
rect 12033 3236 12089 3292
rect 12089 3236 12093 3292
rect 12029 3232 12093 3236
rect 12109 3292 12173 3296
rect 12109 3236 12113 3292
rect 12113 3236 12169 3292
rect 12169 3236 12173 3292
rect 12109 3232 12173 3236
rect 3681 2748 3745 2752
rect 3681 2692 3685 2748
rect 3685 2692 3741 2748
rect 3741 2692 3745 2748
rect 3681 2688 3745 2692
rect 3761 2748 3825 2752
rect 3761 2692 3765 2748
rect 3765 2692 3821 2748
rect 3821 2692 3825 2748
rect 3761 2688 3825 2692
rect 3841 2748 3905 2752
rect 3841 2692 3845 2748
rect 3845 2692 3901 2748
rect 3901 2692 3905 2748
rect 3841 2688 3905 2692
rect 3921 2748 3985 2752
rect 3921 2692 3925 2748
rect 3925 2692 3981 2748
rect 3981 2692 3985 2748
rect 3921 2688 3985 2692
rect 9140 2748 9204 2752
rect 9140 2692 9144 2748
rect 9144 2692 9200 2748
rect 9200 2692 9204 2748
rect 9140 2688 9204 2692
rect 9220 2748 9284 2752
rect 9220 2692 9224 2748
rect 9224 2692 9280 2748
rect 9280 2692 9284 2748
rect 9220 2688 9284 2692
rect 9300 2748 9364 2752
rect 9300 2692 9304 2748
rect 9304 2692 9360 2748
rect 9360 2692 9364 2748
rect 9300 2688 9364 2692
rect 9380 2748 9444 2752
rect 9380 2692 9384 2748
rect 9384 2692 9440 2748
rect 9440 2692 9444 2748
rect 9380 2688 9444 2692
rect 14598 2748 14662 2752
rect 14598 2692 14602 2748
rect 14602 2692 14658 2748
rect 14658 2692 14662 2748
rect 14598 2688 14662 2692
rect 14678 2748 14742 2752
rect 14678 2692 14682 2748
rect 14682 2692 14738 2748
rect 14738 2692 14742 2748
rect 14678 2688 14742 2692
rect 14758 2748 14822 2752
rect 14758 2692 14762 2748
rect 14762 2692 14818 2748
rect 14818 2692 14822 2748
rect 14758 2688 14822 2692
rect 14838 2748 14902 2752
rect 14838 2692 14842 2748
rect 14842 2692 14898 2748
rect 14898 2692 14902 2748
rect 14838 2688 14902 2692
rect 6410 2204 6474 2208
rect 6410 2148 6414 2204
rect 6414 2148 6470 2204
rect 6470 2148 6474 2204
rect 6410 2144 6474 2148
rect 6490 2204 6554 2208
rect 6490 2148 6494 2204
rect 6494 2148 6550 2204
rect 6550 2148 6554 2204
rect 6490 2144 6554 2148
rect 6570 2204 6634 2208
rect 6570 2148 6574 2204
rect 6574 2148 6630 2204
rect 6630 2148 6634 2204
rect 6570 2144 6634 2148
rect 6650 2204 6714 2208
rect 6650 2148 6654 2204
rect 6654 2148 6710 2204
rect 6710 2148 6714 2204
rect 6650 2144 6714 2148
rect 11869 2204 11933 2208
rect 11869 2148 11873 2204
rect 11873 2148 11929 2204
rect 11929 2148 11933 2204
rect 11869 2144 11933 2148
rect 11949 2204 12013 2208
rect 11949 2148 11953 2204
rect 11953 2148 12009 2204
rect 12009 2148 12013 2204
rect 11949 2144 12013 2148
rect 12029 2204 12093 2208
rect 12029 2148 12033 2204
rect 12033 2148 12089 2204
rect 12089 2148 12093 2204
rect 12029 2144 12093 2148
rect 12109 2204 12173 2208
rect 12109 2148 12113 2204
rect 12113 2148 12169 2204
rect 12169 2148 12173 2204
rect 12109 2144 12173 2148
<< metal4 >>
rect 3673 17984 3993 18544
rect 3673 17920 3681 17984
rect 3745 17920 3761 17984
rect 3825 17920 3841 17984
rect 3905 17920 3921 17984
rect 3985 17920 3993 17984
rect 3673 16896 3993 17920
rect 3673 16832 3681 16896
rect 3745 16832 3761 16896
rect 3825 16832 3841 16896
rect 3905 16832 3921 16896
rect 3985 16832 3993 16896
rect 3673 15846 3993 16832
rect 3673 15808 3715 15846
rect 3951 15808 3993 15846
rect 3673 15744 3681 15808
rect 3985 15744 3993 15808
rect 3673 15610 3715 15744
rect 3951 15610 3993 15744
rect 3673 14720 3993 15610
rect 3673 14656 3681 14720
rect 3745 14656 3761 14720
rect 3825 14656 3841 14720
rect 3905 14656 3921 14720
rect 3985 14656 3993 14720
rect 3673 13632 3993 14656
rect 3673 13568 3681 13632
rect 3745 13568 3761 13632
rect 3825 13568 3841 13632
rect 3905 13568 3921 13632
rect 3985 13568 3993 13632
rect 3673 12544 3993 13568
rect 3673 12480 3681 12544
rect 3745 12480 3761 12544
rect 3825 12480 3841 12544
rect 3905 12480 3921 12544
rect 3985 12480 3993 12544
rect 3673 11456 3993 12480
rect 3673 11392 3681 11456
rect 3745 11392 3761 11456
rect 3825 11392 3841 11456
rect 3905 11392 3921 11456
rect 3985 11392 3993 11456
rect 3673 10406 3993 11392
rect 3673 10368 3715 10406
rect 3951 10368 3993 10406
rect 3673 10304 3681 10368
rect 3985 10304 3993 10368
rect 3673 10170 3715 10304
rect 3951 10170 3993 10304
rect 3673 9280 3993 10170
rect 3673 9216 3681 9280
rect 3745 9216 3761 9280
rect 3825 9216 3841 9280
rect 3905 9216 3921 9280
rect 3985 9216 3993 9280
rect 3673 8192 3993 9216
rect 3673 8128 3681 8192
rect 3745 8128 3761 8192
rect 3825 8128 3841 8192
rect 3905 8128 3921 8192
rect 3985 8128 3993 8192
rect 3673 7104 3993 8128
rect 3673 7040 3681 7104
rect 3745 7040 3761 7104
rect 3825 7040 3841 7104
rect 3905 7040 3921 7104
rect 3985 7040 3993 7104
rect 3673 6016 3993 7040
rect 3673 5952 3681 6016
rect 3745 5952 3761 6016
rect 3825 5952 3841 6016
rect 3905 5952 3921 6016
rect 3985 5952 3993 6016
rect 3673 4966 3993 5952
rect 3673 4928 3715 4966
rect 3951 4928 3993 4966
rect 3673 4864 3681 4928
rect 3985 4864 3993 4928
rect 3673 4730 3715 4864
rect 3951 4730 3993 4864
rect 3673 3840 3993 4730
rect 3673 3776 3681 3840
rect 3745 3776 3761 3840
rect 3825 3776 3841 3840
rect 3905 3776 3921 3840
rect 3985 3776 3993 3840
rect 3673 2752 3993 3776
rect 3673 2688 3681 2752
rect 3745 2688 3761 2752
rect 3825 2688 3841 2752
rect 3905 2688 3921 2752
rect 3985 2688 3993 2752
rect 3673 2128 3993 2688
rect 6402 18528 6722 18544
rect 6402 18464 6410 18528
rect 6474 18464 6490 18528
rect 6554 18464 6570 18528
rect 6634 18464 6650 18528
rect 6714 18464 6722 18528
rect 6402 17440 6722 18464
rect 6402 17376 6410 17440
rect 6474 17376 6490 17440
rect 6554 17376 6570 17440
rect 6634 17376 6650 17440
rect 6714 17376 6722 17440
rect 6402 16352 6722 17376
rect 6402 16288 6410 16352
rect 6474 16288 6490 16352
rect 6554 16288 6570 16352
rect 6634 16288 6650 16352
rect 6714 16288 6722 16352
rect 6402 15264 6722 16288
rect 6402 15200 6410 15264
rect 6474 15200 6490 15264
rect 6554 15200 6570 15264
rect 6634 15200 6650 15264
rect 6714 15200 6722 15264
rect 6402 14176 6722 15200
rect 6402 14112 6410 14176
rect 6474 14112 6490 14176
rect 6554 14112 6570 14176
rect 6634 14112 6650 14176
rect 6714 14112 6722 14176
rect 6402 13126 6722 14112
rect 6402 13088 6444 13126
rect 6680 13088 6722 13126
rect 6402 13024 6410 13088
rect 6714 13024 6722 13088
rect 6402 12890 6444 13024
rect 6680 12890 6722 13024
rect 6402 12000 6722 12890
rect 6402 11936 6410 12000
rect 6474 11936 6490 12000
rect 6554 11936 6570 12000
rect 6634 11936 6650 12000
rect 6714 11936 6722 12000
rect 6402 10912 6722 11936
rect 6402 10848 6410 10912
rect 6474 10848 6490 10912
rect 6554 10848 6570 10912
rect 6634 10848 6650 10912
rect 6714 10848 6722 10912
rect 6402 9824 6722 10848
rect 6402 9760 6410 9824
rect 6474 9760 6490 9824
rect 6554 9760 6570 9824
rect 6634 9760 6650 9824
rect 6714 9760 6722 9824
rect 6402 8736 6722 9760
rect 6402 8672 6410 8736
rect 6474 8672 6490 8736
rect 6554 8672 6570 8736
rect 6634 8672 6650 8736
rect 6714 8672 6722 8736
rect 6402 7686 6722 8672
rect 6402 7648 6444 7686
rect 6680 7648 6722 7686
rect 6402 7584 6410 7648
rect 6714 7584 6722 7648
rect 6402 7450 6444 7584
rect 6680 7450 6722 7584
rect 6402 6560 6722 7450
rect 6402 6496 6410 6560
rect 6474 6496 6490 6560
rect 6554 6496 6570 6560
rect 6634 6496 6650 6560
rect 6714 6496 6722 6560
rect 6402 5472 6722 6496
rect 6402 5408 6410 5472
rect 6474 5408 6490 5472
rect 6554 5408 6570 5472
rect 6634 5408 6650 5472
rect 6714 5408 6722 5472
rect 6402 4384 6722 5408
rect 6402 4320 6410 4384
rect 6474 4320 6490 4384
rect 6554 4320 6570 4384
rect 6634 4320 6650 4384
rect 6714 4320 6722 4384
rect 6402 3296 6722 4320
rect 6402 3232 6410 3296
rect 6474 3232 6490 3296
rect 6554 3232 6570 3296
rect 6634 3232 6650 3296
rect 6714 3232 6722 3296
rect 6402 2208 6722 3232
rect 6402 2144 6410 2208
rect 6474 2144 6490 2208
rect 6554 2144 6570 2208
rect 6634 2144 6650 2208
rect 6714 2144 6722 2208
rect 6402 2128 6722 2144
rect 9132 17984 9452 18544
rect 9132 17920 9140 17984
rect 9204 17920 9220 17984
rect 9284 17920 9300 17984
rect 9364 17920 9380 17984
rect 9444 17920 9452 17984
rect 9132 16896 9452 17920
rect 9132 16832 9140 16896
rect 9204 16832 9220 16896
rect 9284 16832 9300 16896
rect 9364 16832 9380 16896
rect 9444 16832 9452 16896
rect 9132 15846 9452 16832
rect 9132 15808 9174 15846
rect 9410 15808 9452 15846
rect 9132 15744 9140 15808
rect 9444 15744 9452 15808
rect 9132 15610 9174 15744
rect 9410 15610 9452 15744
rect 9132 14720 9452 15610
rect 9132 14656 9140 14720
rect 9204 14656 9220 14720
rect 9284 14656 9300 14720
rect 9364 14656 9380 14720
rect 9444 14656 9452 14720
rect 9132 13632 9452 14656
rect 9132 13568 9140 13632
rect 9204 13568 9220 13632
rect 9284 13568 9300 13632
rect 9364 13568 9380 13632
rect 9444 13568 9452 13632
rect 9132 12544 9452 13568
rect 9132 12480 9140 12544
rect 9204 12480 9220 12544
rect 9284 12480 9300 12544
rect 9364 12480 9380 12544
rect 9444 12480 9452 12544
rect 9132 11456 9452 12480
rect 9132 11392 9140 11456
rect 9204 11392 9220 11456
rect 9284 11392 9300 11456
rect 9364 11392 9380 11456
rect 9444 11392 9452 11456
rect 9132 10406 9452 11392
rect 9132 10368 9174 10406
rect 9410 10368 9452 10406
rect 9132 10304 9140 10368
rect 9444 10304 9452 10368
rect 9132 10170 9174 10304
rect 9410 10170 9452 10304
rect 9132 9280 9452 10170
rect 9132 9216 9140 9280
rect 9204 9216 9220 9280
rect 9284 9216 9300 9280
rect 9364 9216 9380 9280
rect 9444 9216 9452 9280
rect 9132 8192 9452 9216
rect 9132 8128 9140 8192
rect 9204 8128 9220 8192
rect 9284 8128 9300 8192
rect 9364 8128 9380 8192
rect 9444 8128 9452 8192
rect 9132 7104 9452 8128
rect 9132 7040 9140 7104
rect 9204 7040 9220 7104
rect 9284 7040 9300 7104
rect 9364 7040 9380 7104
rect 9444 7040 9452 7104
rect 9132 6016 9452 7040
rect 9132 5952 9140 6016
rect 9204 5952 9220 6016
rect 9284 5952 9300 6016
rect 9364 5952 9380 6016
rect 9444 5952 9452 6016
rect 9132 4966 9452 5952
rect 9132 4928 9174 4966
rect 9410 4928 9452 4966
rect 9132 4864 9140 4928
rect 9444 4864 9452 4928
rect 9132 4730 9174 4864
rect 9410 4730 9452 4864
rect 9132 3840 9452 4730
rect 9132 3776 9140 3840
rect 9204 3776 9220 3840
rect 9284 3776 9300 3840
rect 9364 3776 9380 3840
rect 9444 3776 9452 3840
rect 9132 2752 9452 3776
rect 9132 2688 9140 2752
rect 9204 2688 9220 2752
rect 9284 2688 9300 2752
rect 9364 2688 9380 2752
rect 9444 2688 9452 2752
rect 9132 2128 9452 2688
rect 11861 18528 12181 18544
rect 11861 18464 11869 18528
rect 11933 18464 11949 18528
rect 12013 18464 12029 18528
rect 12093 18464 12109 18528
rect 12173 18464 12181 18528
rect 11861 17440 12181 18464
rect 11861 17376 11869 17440
rect 11933 17376 11949 17440
rect 12013 17376 12029 17440
rect 12093 17376 12109 17440
rect 12173 17376 12181 17440
rect 11861 16352 12181 17376
rect 11861 16288 11869 16352
rect 11933 16288 11949 16352
rect 12013 16288 12029 16352
rect 12093 16288 12109 16352
rect 12173 16288 12181 16352
rect 11861 15264 12181 16288
rect 11861 15200 11869 15264
rect 11933 15200 11949 15264
rect 12013 15200 12029 15264
rect 12093 15200 12109 15264
rect 12173 15200 12181 15264
rect 11861 14176 12181 15200
rect 11861 14112 11869 14176
rect 11933 14112 11949 14176
rect 12013 14112 12029 14176
rect 12093 14112 12109 14176
rect 12173 14112 12181 14176
rect 11861 13126 12181 14112
rect 11861 13088 11903 13126
rect 12139 13088 12181 13126
rect 11861 13024 11869 13088
rect 12173 13024 12181 13088
rect 11861 12890 11903 13024
rect 12139 12890 12181 13024
rect 11861 12000 12181 12890
rect 11861 11936 11869 12000
rect 11933 11936 11949 12000
rect 12013 11936 12029 12000
rect 12093 11936 12109 12000
rect 12173 11936 12181 12000
rect 11861 10912 12181 11936
rect 11861 10848 11869 10912
rect 11933 10848 11949 10912
rect 12013 10848 12029 10912
rect 12093 10848 12109 10912
rect 12173 10848 12181 10912
rect 11861 9824 12181 10848
rect 11861 9760 11869 9824
rect 11933 9760 11949 9824
rect 12013 9760 12029 9824
rect 12093 9760 12109 9824
rect 12173 9760 12181 9824
rect 11861 8736 12181 9760
rect 11861 8672 11869 8736
rect 11933 8672 11949 8736
rect 12013 8672 12029 8736
rect 12093 8672 12109 8736
rect 12173 8672 12181 8736
rect 11861 7686 12181 8672
rect 11861 7648 11903 7686
rect 12139 7648 12181 7686
rect 11861 7584 11869 7648
rect 12173 7584 12181 7648
rect 11861 7450 11903 7584
rect 12139 7450 12181 7584
rect 11861 6560 12181 7450
rect 11861 6496 11869 6560
rect 11933 6496 11949 6560
rect 12013 6496 12029 6560
rect 12093 6496 12109 6560
rect 12173 6496 12181 6560
rect 11861 5472 12181 6496
rect 11861 5408 11869 5472
rect 11933 5408 11949 5472
rect 12013 5408 12029 5472
rect 12093 5408 12109 5472
rect 12173 5408 12181 5472
rect 11861 4384 12181 5408
rect 11861 4320 11869 4384
rect 11933 4320 11949 4384
rect 12013 4320 12029 4384
rect 12093 4320 12109 4384
rect 12173 4320 12181 4384
rect 11861 3296 12181 4320
rect 11861 3232 11869 3296
rect 11933 3232 11949 3296
rect 12013 3232 12029 3296
rect 12093 3232 12109 3296
rect 12173 3232 12181 3296
rect 11861 2208 12181 3232
rect 11861 2144 11869 2208
rect 11933 2144 11949 2208
rect 12013 2144 12029 2208
rect 12093 2144 12109 2208
rect 12173 2144 12181 2208
rect 11861 2128 12181 2144
rect 14590 17984 14910 18544
rect 14590 17920 14598 17984
rect 14662 17920 14678 17984
rect 14742 17920 14758 17984
rect 14822 17920 14838 17984
rect 14902 17920 14910 17984
rect 14590 16896 14910 17920
rect 14590 16832 14598 16896
rect 14662 16832 14678 16896
rect 14742 16832 14758 16896
rect 14822 16832 14838 16896
rect 14902 16832 14910 16896
rect 14590 15846 14910 16832
rect 14590 15808 14632 15846
rect 14868 15808 14910 15846
rect 14590 15744 14598 15808
rect 14902 15744 14910 15808
rect 14590 15610 14632 15744
rect 14868 15610 14910 15744
rect 14590 14720 14910 15610
rect 14590 14656 14598 14720
rect 14662 14656 14678 14720
rect 14742 14656 14758 14720
rect 14822 14656 14838 14720
rect 14902 14656 14910 14720
rect 14590 13632 14910 14656
rect 14590 13568 14598 13632
rect 14662 13568 14678 13632
rect 14742 13568 14758 13632
rect 14822 13568 14838 13632
rect 14902 13568 14910 13632
rect 14590 12544 14910 13568
rect 14590 12480 14598 12544
rect 14662 12480 14678 12544
rect 14742 12480 14758 12544
rect 14822 12480 14838 12544
rect 14902 12480 14910 12544
rect 14590 11456 14910 12480
rect 14590 11392 14598 11456
rect 14662 11392 14678 11456
rect 14742 11392 14758 11456
rect 14822 11392 14838 11456
rect 14902 11392 14910 11456
rect 14590 10406 14910 11392
rect 14590 10368 14632 10406
rect 14868 10368 14910 10406
rect 14590 10304 14598 10368
rect 14902 10304 14910 10368
rect 14590 10170 14632 10304
rect 14868 10170 14910 10304
rect 14590 9280 14910 10170
rect 14590 9216 14598 9280
rect 14662 9216 14678 9280
rect 14742 9216 14758 9280
rect 14822 9216 14838 9280
rect 14902 9216 14910 9280
rect 14590 8192 14910 9216
rect 14590 8128 14598 8192
rect 14662 8128 14678 8192
rect 14742 8128 14758 8192
rect 14822 8128 14838 8192
rect 14902 8128 14910 8192
rect 14590 7104 14910 8128
rect 14590 7040 14598 7104
rect 14662 7040 14678 7104
rect 14742 7040 14758 7104
rect 14822 7040 14838 7104
rect 14902 7040 14910 7104
rect 14590 6016 14910 7040
rect 14590 5952 14598 6016
rect 14662 5952 14678 6016
rect 14742 5952 14758 6016
rect 14822 5952 14838 6016
rect 14902 5952 14910 6016
rect 14590 4966 14910 5952
rect 14590 4928 14632 4966
rect 14868 4928 14910 4966
rect 14590 4864 14598 4928
rect 14902 4864 14910 4928
rect 14590 4730 14632 4864
rect 14868 4730 14910 4864
rect 14590 3840 14910 4730
rect 14590 3776 14598 3840
rect 14662 3776 14678 3840
rect 14742 3776 14758 3840
rect 14822 3776 14838 3840
rect 14902 3776 14910 3840
rect 14590 2752 14910 3776
rect 14590 2688 14598 2752
rect 14662 2688 14678 2752
rect 14742 2688 14758 2752
rect 14822 2688 14838 2752
rect 14902 2688 14910 2752
rect 14590 2128 14910 2688
<< via4 >>
rect 3715 15808 3951 15846
rect 3715 15744 3745 15808
rect 3745 15744 3761 15808
rect 3761 15744 3825 15808
rect 3825 15744 3841 15808
rect 3841 15744 3905 15808
rect 3905 15744 3921 15808
rect 3921 15744 3951 15808
rect 3715 15610 3951 15744
rect 3715 10368 3951 10406
rect 3715 10304 3745 10368
rect 3745 10304 3761 10368
rect 3761 10304 3825 10368
rect 3825 10304 3841 10368
rect 3841 10304 3905 10368
rect 3905 10304 3921 10368
rect 3921 10304 3951 10368
rect 3715 10170 3951 10304
rect 3715 4928 3951 4966
rect 3715 4864 3745 4928
rect 3745 4864 3761 4928
rect 3761 4864 3825 4928
rect 3825 4864 3841 4928
rect 3841 4864 3905 4928
rect 3905 4864 3921 4928
rect 3921 4864 3951 4928
rect 3715 4730 3951 4864
rect 6444 13088 6680 13126
rect 6444 13024 6474 13088
rect 6474 13024 6490 13088
rect 6490 13024 6554 13088
rect 6554 13024 6570 13088
rect 6570 13024 6634 13088
rect 6634 13024 6650 13088
rect 6650 13024 6680 13088
rect 6444 12890 6680 13024
rect 6444 7648 6680 7686
rect 6444 7584 6474 7648
rect 6474 7584 6490 7648
rect 6490 7584 6554 7648
rect 6554 7584 6570 7648
rect 6570 7584 6634 7648
rect 6634 7584 6650 7648
rect 6650 7584 6680 7648
rect 6444 7450 6680 7584
rect 9174 15808 9410 15846
rect 9174 15744 9204 15808
rect 9204 15744 9220 15808
rect 9220 15744 9284 15808
rect 9284 15744 9300 15808
rect 9300 15744 9364 15808
rect 9364 15744 9380 15808
rect 9380 15744 9410 15808
rect 9174 15610 9410 15744
rect 9174 10368 9410 10406
rect 9174 10304 9204 10368
rect 9204 10304 9220 10368
rect 9220 10304 9284 10368
rect 9284 10304 9300 10368
rect 9300 10304 9364 10368
rect 9364 10304 9380 10368
rect 9380 10304 9410 10368
rect 9174 10170 9410 10304
rect 9174 4928 9410 4966
rect 9174 4864 9204 4928
rect 9204 4864 9220 4928
rect 9220 4864 9284 4928
rect 9284 4864 9300 4928
rect 9300 4864 9364 4928
rect 9364 4864 9380 4928
rect 9380 4864 9410 4928
rect 9174 4730 9410 4864
rect 11903 13088 12139 13126
rect 11903 13024 11933 13088
rect 11933 13024 11949 13088
rect 11949 13024 12013 13088
rect 12013 13024 12029 13088
rect 12029 13024 12093 13088
rect 12093 13024 12109 13088
rect 12109 13024 12139 13088
rect 11903 12890 12139 13024
rect 11903 7648 12139 7686
rect 11903 7584 11933 7648
rect 11933 7584 11949 7648
rect 11949 7584 12013 7648
rect 12013 7584 12029 7648
rect 12029 7584 12093 7648
rect 12093 7584 12109 7648
rect 12109 7584 12139 7648
rect 11903 7450 12139 7584
rect 14632 15808 14868 15846
rect 14632 15744 14662 15808
rect 14662 15744 14678 15808
rect 14678 15744 14742 15808
rect 14742 15744 14758 15808
rect 14758 15744 14822 15808
rect 14822 15744 14838 15808
rect 14838 15744 14868 15808
rect 14632 15610 14868 15744
rect 14632 10368 14868 10406
rect 14632 10304 14662 10368
rect 14662 10304 14678 10368
rect 14678 10304 14742 10368
rect 14742 10304 14758 10368
rect 14758 10304 14822 10368
rect 14822 10304 14838 10368
rect 14838 10304 14868 10368
rect 14632 10170 14868 10304
rect 14632 4928 14868 4966
rect 14632 4864 14662 4928
rect 14662 4864 14678 4928
rect 14678 4864 14742 4928
rect 14742 4864 14758 4928
rect 14758 4864 14822 4928
rect 14822 4864 14838 4928
rect 14838 4864 14868 4928
rect 14632 4730 14868 4864
<< metal5 >>
rect 1104 15846 17480 15888
rect 1104 15610 3715 15846
rect 3951 15610 9174 15846
rect 9410 15610 14632 15846
rect 14868 15610 17480 15846
rect 1104 15568 17480 15610
rect 1104 13126 17480 13168
rect 1104 12890 6444 13126
rect 6680 12890 11903 13126
rect 12139 12890 17480 13126
rect 1104 12848 17480 12890
rect 1104 10406 17480 10448
rect 1104 10170 3715 10406
rect 3951 10170 9174 10406
rect 9410 10170 14632 10406
rect 14868 10170 17480 10406
rect 1104 10128 17480 10170
rect 1104 7686 17480 7728
rect 1104 7450 6444 7686
rect 6680 7450 11903 7686
rect 12139 7450 17480 7686
rect 1104 7408 17480 7450
rect 1104 4966 17480 5008
rect 1104 4730 3715 4966
rect 3951 4730 9174 4966
rect 9410 4730 14632 4966
rect 14868 4730 17480 4966
rect 1104 4688 17480 4730
use sky130_fd_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1631199322
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1631199322
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1631199322
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1631199322
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1631199322
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1631199322
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1631199322
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1631199322
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1631199322
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1631199322
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45
timestamp 1631199322
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1631199322
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1631199322
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1631199322
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1631199322
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1631199322
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1631199322
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1631199322
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1631199322
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 6808 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _43_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 6808 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1631199322
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1631199322
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1631199322
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _30_
timestamp 1631199322
transform -1 0 8464 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1631199322
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1631199322
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _44_
timestamp 1631199322
transform 1 0 9016 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_sclk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 9200 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1631199322
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1631199322
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1631199322
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1631199322
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1631199322
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1631199322
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _25_
timestamp 1631199322
transform 1 0 12236 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _46_
timestamp 1631199322
transform 1 0 11960 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_138
timestamp 1631199322
transform 1 0 13800 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1631199322
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1631199322
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1631199322
transform -1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1631199322
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _28_
timestamp 1631199322
transform -1 0 14720 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_1_150
timestamp 1631199322
transform 1 0 14904 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1631199322
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1631199322
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1631199322
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1631199322
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1631199322
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1631199322
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1631199322
transform -1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1631199322
transform -1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1631199322
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1631199322
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1631199322
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1631199322
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1631199322
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1631199322
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1631199322
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1631199322
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1631199322
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1631199322
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1631199322
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_sclk
timestamp 1631199322
transform -1 0 7084 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1631199322
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1631199322
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1631199322
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1631199322
transform -1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_95
timestamp 1631199322
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1631199322
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1631199322
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _45_
timestamp 1631199322
transform 1 0 10212 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1631199322
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1631199322
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _22_
timestamp 1631199322
transform 1 0 12604 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_119
timestamp 1631199322
transform 1 0 12052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_145
timestamp 1631199322
transform 1 0 14444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1631199322
transform -1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1631199322
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1631199322
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_157
timestamp 1631199322
transform 1 0 15548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1631199322
transform -1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_169
timestamp 1631199322
transform 1 0 16652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1631199322
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1631199322
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1631199322
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1631199322
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1631199322
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1631199322
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1631199322
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1631199322
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1631199322
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1631199322
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _34_
timestamp 1631199322
transform 1 0 6808 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1631199322
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1631199322
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _36_
timestamp 1631199322
transform 1 0 8464 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1631199322
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1631199322
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_87
timestamp 1631199322
transform 1 0 9108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 10396 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1631199322
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_116
timestamp 1631199322
transform 1 0 11776 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1631199322
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _47_
timestamp 1631199322
transform 1 0 12512 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1631199322
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1631199322
transform 1 0 14352 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1631199322
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1631199322
transform -1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1631199322
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1631199322
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1631199322
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1631199322
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1631199322
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1631199322
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1631199322
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1631199322
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1631199322
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1631199322
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1631199322
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _42_
timestamp 1631199322
transform 1 0 6440 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1631199322
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1631199322
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1631199322
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_sclk
timestamp 1631199322
transform 1 0 9568 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1631199322
transform 1 0 8924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp 1631199322
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1631199322
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _24_
timestamp 1631199322
transform -1 0 13156 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1631199322
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1631199322
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1631199322
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1631199322
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1631199322
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_148
timestamp 1631199322
transform 1 0 14720 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_160
timestamp 1631199322
transform 1 0 15824 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_172
timestamp 1631199322
transform 1 0 16928 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1631199322
transform -1 0 17480 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1631199322
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1631199322
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1631199322
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1631199322
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1631199322
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1631199322
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1631199322
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1631199322
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1631199322
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1631199322
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _41_
timestamp 1631199322
transform -1 0 8832 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_5_84
timestamp 1631199322
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _40_
timestamp 1631199322
transform -1 0 11040 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1631199322
transform 1 0 12420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1631199322
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1631199322
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _27_
timestamp 1631199322
transform -1 0 12420 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1631199322
transform 1 0 13524 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1631199322
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_159
timestamp 1631199322
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1631199322
transform -1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1631199322
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1631199322
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_169
timestamp 1631199322
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1631199322
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1631199322
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1631199322
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1631199322
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1631199322
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1631199322
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1631199322
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1631199322
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1631199322
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1631199322
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1631199322
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1631199322
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1631199322
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1631199322
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1631199322
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1631199322
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1631199322
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1631199322
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1631199322
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1631199322
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1631199322
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1631199322
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1631199322
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1631199322
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1631199322
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _38_
timestamp 1631199322
transform 1 0 10396 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1631199322
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_94
timestamp 1631199322
transform 1 0 9752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1631199322
transform 1 0 9476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_120
timestamp 1631199322
transform 1 0 12144 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1631199322
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1631199322
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_116
timestamp 1631199322
transform 1 0 11776 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1631199322
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_108
timestamp 1631199322
transform 1 0 11040 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1631199322
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1631199322
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1631199322
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1631199322
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1631199322
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_132
timestamp 1631199322
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1631199322
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1631199322
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1631199322
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_165
timestamp 1631199322
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1631199322
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1631199322
transform -1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1631199322
transform -1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1631199322
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1631199322
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_169
timestamp 1631199322
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_173 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform 1 0 17020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1631199322
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1631199322
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1631199322
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1631199322
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1631199322
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1631199322
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1631199322
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1631199322
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1631199322
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1631199322
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1631199322
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1631199322
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1631199322
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1631199322
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1631199322
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1631199322
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1631199322
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1631199322
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1631199322
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1631199322
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1631199322
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_165
timestamp 1631199322
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1631199322
transform -1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_173
timestamp 1631199322
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1631199322
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1631199322
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1631199322
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1631199322
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1631199322
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1631199322
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1631199322
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1631199322
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1631199322
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1631199322
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1631199322
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1631199322
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1631199322
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1631199322
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1631199322
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1631199322
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1631199322
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1631199322
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1631199322
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1631199322
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1631199322
transform -1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1631199322
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1631199322
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1631199322
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1631199322
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1631199322
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1631199322
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1631199322
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1631199322
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1631199322
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1631199322
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1631199322
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1631199322
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1631199322
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1631199322
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1631199322
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1631199322
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1631199322
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1631199322
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1631199322
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1631199322
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1631199322
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1631199322
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1631199322
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1631199322
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1631199322
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1631199322
transform -1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1631199322
transform 1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1631199322
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1631199322
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1631199322
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1631199322
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1631199322
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1631199322
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1631199322
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1631199322
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1631199322
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1631199322
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1631199322
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1631199322
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1631199322
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1631199322
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1631199322
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1631199322
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1631199322
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1631199322
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1631199322
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1631199322
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1631199322
transform -1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1631199322
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1631199322
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_169
timestamp 1631199322
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1631199322
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1631199322
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1631199322
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1631199322
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1631199322
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1631199322
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1631199322
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1631199322
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1631199322
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1631199322
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1631199322
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1631199322
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1631199322
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1631199322
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1631199322
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1631199322
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1631199322
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1631199322
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1631199322
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1631199322
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1631199322
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp 1631199322
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1631199322
transform -1 0 17480 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1631199322
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1631199322
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1631199322
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1631199322
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1631199322
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1631199322
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1631199322
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1631199322
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1631199322
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1631199322
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1631199322
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1631199322
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1631199322
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1631199322
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1631199322
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1631199322
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1631199322
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1631199322
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1631199322
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1631199322
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1631199322
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1631199322
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1631199322
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1631199322
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1631199322
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1631199322
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1631199322
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1631199322
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1631199322
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1631199322
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1631199322
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1631199322
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1631199322
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1631199322
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1631199322
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1631199322
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1631199322
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1631199322
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1631199322
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1631199322
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1631199322
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_165
timestamp 1631199322
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1631199322
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1631199322
transform -1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1631199322
transform -1 0 17480 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1631199322
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1631199322
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1631199322
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_173
timestamp 1631199322
transform 1 0 17020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1631199322
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1631199322
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1631199322
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1631199322
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1631199322
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1631199322
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1631199322
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1631199322
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1631199322
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1631199322
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1631199322
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1631199322
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1631199322
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1631199322
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1631199322
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1631199322
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1631199322
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1631199322
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1631199322
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1631199322
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1631199322
transform -1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1631199322
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1631199322
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1631199322
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1631199322
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1631199322
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1631199322
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1631199322
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1631199322
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1631199322
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1631199322
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1631199322
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1631199322
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1631199322
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1631199322
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1631199322
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1631199322
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1631199322
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1631199322
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1631199322
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1631199322
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1631199322
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1631199322
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1631199322
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1631199322
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1631199322
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1631199322
transform -1 0 17480 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1631199322
transform 1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1631199322
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1631199322
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1631199322
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1631199322
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1631199322
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1631199322
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1631199322
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1631199322
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1631199322
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1631199322
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1631199322
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1631199322
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1631199322
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1631199322
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1631199322
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1631199322
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1631199322
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1631199322
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1631199322
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1631199322
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1631199322
transform -1 0 17480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1631199322
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1631199322
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1631199322
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1631199322
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1631199322
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1631199322
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1631199322
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1631199322
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1631199322
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1631199322
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1631199322
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1631199322
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1631199322
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1631199322
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1631199322
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1631199322
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1631199322
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1631199322
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1631199322
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1631199322
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1631199322
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1631199322
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1631199322
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1631199322
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_165
timestamp 1631199322
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1631199322
transform -1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp 1631199322
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1631199322
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1631199322
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1631199322
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1631199322
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1631199322
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1631199322
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1631199322
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1631199322
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1631199322
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1631199322
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1631199322
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1631199322
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1631199322
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1631199322
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1631199322
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1631199322
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1631199322
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1631199322
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1631199322
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1631199322
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1631199322
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1631199322
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1631199322
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1631199322
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1631199322
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1631199322
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1631199322
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1631199322
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1631199322
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1631199322
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1631199322
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1631199322
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1631199322
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1631199322
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1631199322
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1631199322
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1631199322
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1631199322
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1631199322
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1631199322
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_165
timestamp 1631199322
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1631199322
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1631199322
transform -1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1631199322
transform -1 0 17480 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1631199322
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1631199322
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1631199322
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_173
timestamp 1631199322
transform 1 0 17020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1631199322
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1631199322
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1631199322
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1631199322
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1631199322
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1631199322
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1631199322
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1631199322
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1631199322
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1631199322
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1631199322
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1631199322
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1631199322
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1631199322
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1631199322
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1631199322
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1631199322
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1631199322
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1631199322
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1631199322
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1631199322
transform -1 0 17480 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1631199322
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1631199322
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1631199322
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1631199322
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1631199322
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1631199322
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1631199322
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1631199322
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1631199322
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1631199322
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1631199322
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1631199322
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1631199322
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1631199322
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1631199322
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1631199322
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1631199322
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1631199322
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1631199322
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1631199322
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1631199322
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1631199322
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1631199322
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1631199322
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_165
timestamp 1631199322
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1631199322
transform -1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_173
timestamp 1631199322
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1631199322
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1631199322
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1631199322
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1631199322
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1631199322
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1631199322
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1631199322
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1631199322
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1631199322
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1631199322
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1631199322
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1631199322
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1631199322
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1631199322
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1631199322
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1631199322
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1631199322
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1631199322
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1631199322
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1631199322
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1631199322
transform -1 0 17480 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1631199322
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1631199322
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 1631199322
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1631199322
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1631199322
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1631199322
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1631199322
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1631199322
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1631199322
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1631199322
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1631199322
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1631199322
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1631199322
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1631199322
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1631199322
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1631199322
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1631199322
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1631199322
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1631199322
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1631199322
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1631199322
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1631199322
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1631199322
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1631199322
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_165
timestamp 1631199322
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1631199322
transform -1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1631199322
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1631199322
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1631199322
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1631199322
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1631199322
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1631199322
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1631199322
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1631199322
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1631199322
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1631199322
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1631199322
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1631199322
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1631199322
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1631199322
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1631199322
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1631199322
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1631199322
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1631199322
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1631199322
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1631199322
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1631199322
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1631199322
transform -1 0 17480 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1631199322
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1631199322
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1631199322
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1631199322
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1631199322
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1631199322
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1631199322
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1631199322
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1631199322
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1631199322
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1631199322
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1631199322
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1631199322
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1631199322
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1631199322
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1631199322
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1631199322
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1631199322
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1631199322
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1631199322
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1631199322
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1631199322
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1631199322
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1631199322
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1631199322
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1631199322
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1631199322
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1631199322
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1631199322
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1631199322
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1631199322
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1631199322
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1631199322
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1631199322
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1631199322
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1631199322
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1631199322
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1631199322
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1631199322
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1631199322
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1631199322
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1631199322
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1631199322
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_165
timestamp 1631199322
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1631199322
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1631199322
transform -1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1631199322
transform -1 0 17480 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1631199322
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1631199322
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1631199322
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1631199322
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1631199322
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1631199322
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1631199322
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1631199322
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1631199322
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1631199322
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1631199322
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1631199322
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1631199322
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1631199322
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1631199322
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1631199322
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1631199322
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1631199322
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1631199322
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1631199322
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1631199322
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1631199322
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1631199322
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1631199322
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_161
timestamp 1631199322
transform 1 0 15916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1631199322
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_157
timestamp 1631199322
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _23_
timestamp 1631199322
transform -1 0 15916 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1631199322
transform -1 0 17480 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1631199322
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_11
timestamp 1631199322
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1631199322
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1631199322
transform 1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_18
timestamp 1631199322
transform 1 0 2760 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1631199322
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1631199322
transform 1 0 3772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_41
timestamp 1631199322
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1631199322
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1631199322
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1631199322
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1631199322
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1631199322
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1631199322
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_81
timestamp 1631199322
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_85
timestamp 1631199322
transform 1 0 8924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_97
timestamp 1631199322
transform 1 0 10028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1631199322
transform 1 0 8832 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_118
timestamp 1631199322
transform 1 0 11960 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1631199322
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1631199322
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1631199322
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631199322
transform -1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1631199322
transform 1 0 14076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_130
timestamp 1631199322
transform 1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1631199322
transform 1 0 13984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1631199322
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1631199322
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_153
timestamp 1631199322
transform 1 0 15180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1631199322
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1631199322
transform -1 0 17480 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1631199322
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1631199322
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
<< labels >>
rlabel metal5 s 1104 7408 17480 7728 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 4688 17480 5008 6 VPWR
port 1 nsew power input
rlabel metal2 s 1122 0 1178 800 6 data[0]
port 2 nsew signal tristate
rlabel metal2 s 3422 0 3478 800 6 data[1]
port 3 nsew signal tristate
rlabel metal2 s 5722 0 5778 800 6 data[2]
port 4 nsew signal tristate
rlabel metal2 s 8022 0 8078 800 6 data[3]
port 5 nsew signal tristate
rlabel metal2 s 10414 0 10470 800 6 data[4]
port 6 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 data[5]
port 7 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 data[6]
port 8 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 data[7]
port 9 nsew signal tristate
rlabel metal2 s 16210 19931 16266 20731 6 reset
port 10 nsew signal input
rlabel metal2 s 6918 19931 6974 20731 6 sclk
port 11 nsew signal input
rlabel metal2 s 11610 19931 11666 20731 6 sdi
port 12 nsew signal input
rlabel metal2 s 2318 19931 2374 20731 6 ss
port 13 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 18587 20731
<< end >>
