*TB CMRR OTA BUFFERED

.include ./ota.spice

X1	IN1	IN1	VD	VS	A	OUT ota

CL	OUT	0	4p

Ibias A 0 5.53u

VDD VD 0 1.8
VSS VS 0 -1.8

*CMRR

*Modo comum
VIN1 IN1 0 DC 0 AC 1

* cmd 	step	stop
.ac	dec	2000	1	110Meg

.end

.control

destroy all
run

*CMRR
plot db(OUT) 

.endc
