*tb-digpot
.include ./digpot.spice
.include ../minimal_libs/sky130_libs/sky130_lib.spice

Xdp	n8	0	vdd	vss	c7 c6 c5 c4 c3 c2 c1 c0 digpot

Vdd	vdd	0	1.8
Vss	vss	0	0

V8	n8	0	1.8

Vc7	c7	0	pulse(1.8 0 0 0 0 640m 1280m)
Vc6	c6	0	pulse(1.8 0 0 0 0 320m 640m)
Vc5	c5	0	pulse(1.8 0 0 0 0 160m 320m)
Vc4	c4	0	pulse(1.8 0 0 0 0 80m 160m)
Vc3	c3	0	pulse(1.8 0 0 0 0 40m 80m)
Vc2	c2	0	pulse(1.8 0 0 0 0 20m 40m)
Vc1	c1	0	pulse(1.8 0 0 0 0 10m 20m)
Vc0	c0	0	pulse(1.8 0 0 0 0 5m 10m)

.end

.control

run

tran 1m 1280m 5m
let Rf=abs(n8/i(V8))
plot Rf

plot c0 c1+2 c2+4 c3+6 c4+8 c6+10 c7+12

.endc
