** transmission gate **

.include ../minimal_libs/sky130_libs/sky130_lib.spice

.subckt	tg	ctrl	a	b	vdd	vss

*lbl	drain	gate	source	bulk	model			length	width
xm1	b	nctrl	a	vss	sky130_fd_pr__nfet_01v8	L=0.15u	W=1u
xm2	a	ctrl	b	vdd	sky130_fd_pr__pfet_01v8	L=0.15u	W=3u
xm3	nctrl	ctrl	vdd	vdd	sky130_fd_pr__pfet_01v8	L=0.15u	W=3u
xm4	nctrl	ctrl	vss	vss	sky130_fd_pr__nfet_01v8	L=0.15u	W=1u

.ends
