magic
tech sky130A
magscale 1 2
timestamp 1634750299
<< nwell >>
rect 2660 7690 2860 7810
rect 3880 7690 4080 7810
rect 4150 7710 4310 7770
rect 4410 7710 4570 7770
rect 4670 7710 4830 7770
rect 4930 7710 5090 7770
rect 6140 7710 6300 7770
rect 1320 6520 1500 6740
<< pmos >>
rect 2660 7779 2856 7810
rect 3880 7779 4076 7810
<< pdiff >>
rect 2856 7779 2860 7810
rect 4076 7779 4080 7810
<< poly >>
rect 2660 7732 2856 7779
rect 2660 7698 2672 7732
rect 2840 7698 2856 7732
rect 2660 7690 2856 7698
rect 3880 7732 4076 7779
rect 3880 7698 3892 7732
rect 4060 7698 4076 7732
rect 4150 7710 4310 7770
rect 4410 7710 4570 7770
rect 4670 7710 4830 7770
rect 4930 7710 5090 7770
rect 6140 7710 6300 7770
rect 3880 7690 4076 7698
<< polycont >>
rect 2672 7698 2840 7732
rect 3892 7698 4060 7732
<< locali >>
rect 2660 7698 2672 7732
rect 2840 7698 2856 7732
rect 3880 7698 3892 7732
rect 4060 7698 4076 7732
<< viali >>
rect 2672 7698 2840 7732
rect 3892 7698 4060 7732
<< metal1 >>
rect -480 9660 -280 9860
rect 0 9660 200 9860
rect 1120 9660 1320 9860
rect -1120 7520 -700 7560
rect -1120 7380 -880 7520
rect -740 7380 -700 7520
rect -1120 7340 -700 7380
rect -500 5910 -250 9660
rect -20 6190 230 9660
rect 1060 9440 1400 9660
rect 1060 9080 6480 9440
rect 1060 8940 1400 9080
rect 2340 8940 2600 9080
rect 3550 8940 3830 9080
rect 5780 8940 6020 9080
rect 1060 8460 1580 8940
rect 1800 8140 2180 8600
rect 2340 8460 2640 8940
rect 3550 8700 5160 8940
rect 2860 8140 3340 8600
rect 3550 8470 3830 8700
rect 5780 8460 6120 8940
rect 1600 7770 1790 7810
rect 1600 7710 1610 7770
rect 1770 7710 1790 7770
rect 1600 7690 1790 7710
rect 1960 7560 2180 8140
rect 2660 7770 2850 7810
rect 2660 7710 2670 7770
rect 2830 7738 2850 7770
rect 2830 7732 2852 7738
rect 2660 7698 2672 7710
rect 2840 7698 2852 7732
rect 2660 7692 2852 7698
rect 2660 7690 2850 7692
rect 440 7520 2180 7560
rect 440 7380 500 7520
rect 720 7380 2180 7520
rect 3080 7500 3340 8140
rect 4080 8130 5450 8370
rect 6330 8130 6760 8600
rect 3880 7770 4070 7810
rect 3880 7710 3890 7770
rect 4050 7738 4070 7770
rect 4130 7770 4340 7790
rect 4050 7732 4072 7738
rect 3880 7698 3892 7710
rect 4060 7698 4072 7732
rect 3880 7692 4072 7698
rect 4130 7710 4150 7770
rect 4310 7710 4340 7770
rect 3880 7690 4070 7692
rect 4130 7680 4340 7710
rect 4390 7770 4590 7780
rect 4390 7710 4410 7770
rect 4570 7710 4590 7770
rect 4390 7680 4590 7710
rect 4650 7770 4850 7780
rect 4650 7710 4670 7770
rect 4830 7710 4850 7770
rect 4650 7680 4850 7710
rect 4910 7770 5110 7780
rect 4910 7710 4930 7770
rect 5090 7710 5110 7770
rect 4910 7680 5110 7710
rect 440 7340 2180 7380
rect 2260 7340 3340 7500
rect 1460 7240 2140 7250
rect 2260 7240 3000 7340
rect 5270 7290 5450 8130
rect 6120 7770 6320 7780
rect 6120 7710 6140 7770
rect 6300 7710 6320 7770
rect 6120 7680 6320 7710
rect 1460 7080 3000 7240
rect 1460 7070 2540 7080
rect 2850 7070 3000 7080
rect 1900 6900 2540 7070
rect 4180 7020 5450 7290
rect -20 6080 40 6190
rect 170 6080 230 6190
rect -20 6050 230 6080
rect 1300 6520 1580 6740
rect 1800 6680 2640 6900
rect 2860 6520 3280 6740
rect 4970 6690 5450 7020
rect 6500 7170 6760 8130
rect 6500 6970 6960 7170
rect 6500 6780 6760 6970
rect 4970 6640 5340 6690
rect -500 5800 -450 5910
rect -320 5800 -250 5910
rect -500 5760 -250 5800
rect 1300 5820 1440 6520
rect 1600 6320 1790 6340
rect 1600 6260 1620 6320
rect 1780 6260 1790 6320
rect 1600 6250 1790 6260
rect 2660 6320 2850 6340
rect 2660 6260 2670 6320
rect 2830 6260 2850 6320
rect 2660 6240 2850 6260
rect 3020 6010 3280 6520
rect 4520 6490 5020 6640
rect 5320 6490 5340 6640
rect 5980 6540 6760 6780
rect 4520 6440 5340 6490
rect 5380 6430 6320 6490
rect 5380 6400 6310 6430
rect 5380 6240 5600 6400
rect 6500 6380 6760 6540
rect 4270 6050 5600 6240
rect 4970 6010 5210 6050
rect 3020 5860 5210 6010
rect 1300 5620 2860 5820
rect 1300 5360 1440 5620
rect 1580 5400 1780 5620
rect 2660 5400 2860 5620
rect 3020 5400 3280 5860
rect 3020 5360 3120 5400
rect 1300 5260 1580 5360
rect 1780 5190 2650 5350
rect 2860 5290 3120 5360
rect 3270 5290 3280 5400
rect 2860 5260 3280 5290
rect 1940 5060 2490 5190
rect 4970 5060 5210 5860
rect 5640 5570 6110 6030
rect 6330 5900 6760 6380
rect 5640 5060 5920 5570
rect 1440 4990 6760 5060
rect 1440 4790 6960 4990
rect 1440 4720 6760 4790
<< via1 >>
rect -880 7380 -740 7520
rect 1610 7710 1770 7770
rect 2670 7732 2830 7770
rect 2670 7710 2672 7732
rect 2672 7710 2830 7732
rect 500 7380 720 7520
rect 3890 7732 4050 7770
rect 3890 7710 3892 7732
rect 3892 7710 4050 7732
rect 4150 7710 4310 7770
rect 4410 7710 4570 7770
rect 4670 7710 4830 7770
rect 4930 7710 5090 7770
rect 6140 7710 6300 7770
rect 40 6080 170 6190
rect -450 5800 -320 5910
rect 1620 6260 1780 6320
rect 2670 6260 2830 6320
rect 5020 6490 5320 6640
rect 3120 5290 3270 5400
<< metal2 >>
rect 1540 7770 6330 7830
rect 1540 7710 1610 7770
rect 1770 7710 2670 7770
rect 2830 7710 3890 7770
rect 4050 7710 4150 7770
rect 4310 7710 4410 7770
rect 4570 7710 4670 7770
rect 4830 7710 4930 7770
rect 5090 7710 6140 7770
rect 6300 7710 6330 7770
rect 1540 7680 6330 7710
rect -920 7520 780 7560
rect -920 7380 -880 7520
rect -740 7380 500 7520
rect 720 7380 780 7520
rect -920 7340 780 7380
rect 4990 6640 5350 6700
rect 4990 6490 5020 6640
rect 5320 6490 5350 6640
rect 1600 6320 1810 6340
rect 1600 6260 1620 6320
rect 1780 6260 1810 6320
rect 1600 6230 1810 6260
rect -20 6190 1810 6230
rect -20 6080 40 6190
rect 170 6080 1810 6190
rect -20 6050 1810 6080
rect 2650 6320 2860 6340
rect 2650 6260 2670 6320
rect 2830 6260 2860 6320
rect 2650 5940 2860 6260
rect -500 5910 2860 5940
rect -500 5800 -450 5910
rect -320 5800 2860 5910
rect -500 5760 2860 5800
rect 3060 5400 3310 5440
rect 3060 5290 3120 5400
rect 3270 5290 3310 5400
rect 3060 4520 3310 5290
rect 3060 4410 3110 4520
rect 3260 4410 3310 4520
rect 3060 4360 3310 4410
rect 4990 4580 5350 6490
rect 4990 4340 6500 4580
rect 6180 4180 6500 4340
rect 6180 4010 6240 4180
rect 6430 4010 6500 4180
rect 6180 3920 6500 4010
<< via2 >>
rect 3110 4410 3260 4520
rect 6240 4010 6430 4180
<< metal3 >>
rect 3060 4520 3310 4580
rect 3060 4410 3110 4520
rect 3260 4410 3310 4520
rect 3060 3990 3310 4410
rect 6180 4180 6500 4300
rect 6180 4010 6240 4180
rect 6430 4010 6500 4180
rect 6180 3920 6500 4010
<< via3 >>
rect 6240 4010 6430 4180
<< metal4 >>
rect 5940 4180 6490 4290
rect 5940 4010 6240 4180
rect 6430 4010 6490 4180
rect 5940 3930 6490 4010
use sky130_fd_pr__cap_mim_m3_1_UYJ6HG  XCC
timestamp 1634487483
transform 1 0 3682 0 1 2002
box -2352 -2302 2351 2302
use sky130_fd_pr__pfet_01v8_5LYT2L  XM2
timestamp 1634510737
transform 1 0 2756 0 1 6632
box -296 -512 296 512
use sky130_fd_pr__nfet_01v8_WJ5JTF  XM4
timestamp 1634510737
transform -1 0 2756 0 1 5276
box -296 -296 296 296
use sky130_fd_pr__pfet_01v8_YRRRD6  XM1
timestamp 1634510737
transform -1 0 1696 0 1 6632
box -296 -512 296 512
use sky130_fd_pr__nfet_01v8_NYLAJZ  XM3
timestamp 1634510737
transform 1 0 1676 0 1 5276
box -296 -296 296 296
use sky130_fd_pr__nfet_01v8_GVU33C  XM7
timestamp 1634510737
transform -1 0 4545 0 -1 6461
box -425 -641 425 641
use sky130_fd_pr__pfet_01v8_UPMF5R  XM9
timestamp 1634510737
transform -1 0 6216 0 1 5804
box -296 -804 296 804
use sky130_fd_pr__pfet_01v8_W5QVET  XM6
timestamp 1634510737
transform 1 0 2756 0 1 8364
box -296 -804 296 804
use sky130_fd_pr__pfet_01v8_W5QVET  XM5
timestamp 1634510737
transform 1 0 1696 0 1 8364
box -296 -804 296 804
use sky130_fd_pr__pfet_01v8_W7P4FT  XM8
timestamp 1634510737
transform 1 0 4492 0 1 8365
box -812 -805 812 805
use sky130_fd_pr__pfet_01v8_W5QVET  XM10
timestamp 1634510737
transform 1 0 6216 0 1 8364
box -296 -804 296 804
<< labels >>
flabel metal1 1120 9660 1320 9860 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 -480 9660 -280 9860 0 FreeSans 256 0 0 0 in1
port 3 nsew
flabel metal1 0 9660 200 9860 0 FreeSans 256 0 0 0 in2
port 4 nsew
flabel metal1 6760 4790 6960 4990 0 FreeSans 256 0 0 0 vs
port 1 nsew
flabel metal1 6760 6970 6960 7170 0 FreeSans 256 0 0 0 out
port 5 nsew
flabel metal1 -1120 7360 -920 7560 0 FreeSans 256 0 0 0 ib
port 2 nsew
<< end >>
