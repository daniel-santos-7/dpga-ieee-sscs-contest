
.include	../minimal_libs/pshort.lib
.include	../minimal_libs/nshort.lib
.include	./tg.spice

.subckt	digpot	n0	n8	vdd	vss	c7 c6 c5 c4 c3 c2 c1 c0	Rn=850

Xtg7	c7	n8	n7	vdd	vss	tg
Xtg6	c6	n7	n6	vdd	vss	tg
Xtg5	c5	n6	n5	vdd	vss	tg
Xtg4	c4	n5	n4	vdd	vss	tg
Xtg3	c3	n4	n3	vdd	vss	tg
Xtg2	c2	n3	n2	vdd	vss	tg
Xtg1	c1	n2	n1	vdd	vss	tg
Xtg0	c0	n1	n0	vdd	vss	tg

R7	n8	n7	{128*Rn}
R6	n7	n6	{64*Rn}
R5	n6	n5	{32*Rn}
R4	n5	n4	{16*Rn}
R3	n4	n3	{8*Rn}
R2	n3	n2	{4*Rn}
R1	n2	n1	{2*Rn}
R0	n1	n0	{Rn}

.ends

